magic
tech sky130A
magscale 1 2
timestamp 1698770908
<< metal1 >>
rect 338298 85212 338304 85264
rect 338356 85252 338362 85264
rect 338666 85252 338672 85264
rect 338356 85224 338672 85252
rect 338356 85212 338362 85224
rect 338666 85212 338672 85224
rect 338724 85212 338730 85264
rect 337378 80248 337384 80300
rect 337436 80248 337442 80300
rect 337396 80096 337424 80248
rect 336550 80044 336556 80096
rect 336608 80084 336614 80096
rect 336734 80084 336740 80096
rect 336608 80056 336740 80084
rect 336608 80044 336614 80056
rect 336734 80044 336740 80056
rect 336792 80044 336798 80096
rect 337378 80044 337384 80096
rect 337436 80044 337442 80096
rect 81756 79908 81762 79960
rect 81814 79948 81820 79960
rect 398098 79948 398104 79960
rect 81814 79920 398104 79948
rect 81814 79908 81820 79920
rect 398098 79908 398104 79920
rect 398156 79908 398162 79960
rect 338850 79432 338856 79484
rect 338908 79432 338914 79484
rect 338868 79280 338896 79432
rect 338850 79228 338856 79280
rect 338908 79228 338914 79280
rect 124122 78616 124128 78668
rect 124180 78656 124186 78668
rect 173986 78656 173992 78668
rect 124180 78628 173992 78656
rect 124180 78616 124186 78628
rect 173986 78616 173992 78628
rect 174044 78616 174050 78668
rect 178034 78616 178040 78668
rect 178092 78656 178098 78668
rect 329466 78656 329472 78668
rect 178092 78628 329472 78656
rect 178092 78616 178098 78628
rect 329466 78616 329472 78628
rect 329524 78616 329530 78668
rect 118694 78548 118700 78600
rect 118752 78588 118758 78600
rect 152090 78588 152096 78600
rect 118752 78560 152096 78588
rect 118752 78548 118758 78560
rect 152090 78548 152096 78560
rect 152148 78548 152154 78600
rect 117222 78480 117228 78532
rect 117280 78520 117286 78532
rect 142706 78520 142712 78532
rect 117280 78492 142712 78520
rect 117280 78480 117286 78492
rect 142706 78480 142712 78492
rect 142764 78480 142770 78532
rect 320818 78140 320824 78192
rect 320876 78180 320882 78192
rect 400950 78180 400956 78192
rect 320876 78152 400956 78180
rect 320876 78140 320882 78152
rect 400950 78140 400956 78152
rect 401008 78140 401014 78192
rect 305638 78072 305644 78124
rect 305696 78112 305702 78124
rect 408770 78112 408776 78124
rect 305696 78084 408776 78112
rect 305696 78072 305702 78084
rect 408770 78072 408776 78084
rect 408828 78072 408834 78124
rect 174538 78004 174544 78056
rect 174596 78044 174602 78056
rect 302418 78044 302424 78056
rect 174596 78016 302424 78044
rect 174596 78004 174602 78016
rect 302418 78004 302424 78016
rect 302476 78004 302482 78056
rect 307018 78004 307024 78056
rect 307076 78044 307082 78056
rect 411898 78044 411904 78056
rect 307076 78016 411904 78044
rect 307076 78004 307082 78016
rect 411898 78004 411904 78016
rect 411956 78004 411962 78056
rect 181438 77936 181444 77988
rect 181496 77976 181502 77988
rect 333974 77976 333980 77988
rect 181496 77948 333980 77976
rect 181496 77936 181502 77948
rect 333974 77936 333980 77948
rect 334032 77936 334038 77988
rect 144914 77800 144920 77852
rect 144972 77840 144978 77852
rect 146018 77840 146024 77852
rect 144972 77812 146024 77840
rect 144972 77800 144978 77812
rect 146018 77800 146024 77812
rect 146076 77800 146082 77852
rect 75822 12384 75828 12436
rect 75880 12424 75886 12436
rect 191282 12424 191288 12436
rect 75880 12396 191288 12424
rect 75880 12384 75886 12396
rect 191282 12384 191288 12396
rect 191340 12384 191346 12436
rect 78582 12316 78588 12368
rect 78640 12356 78646 12368
rect 191190 12356 191196 12368
rect 78640 12328 191196 12356
rect 78640 12316 78646 12328
rect 191190 12316 191196 12328
rect 191248 12316 191254 12368
rect 88242 10956 88248 11008
rect 88300 10996 88306 11008
rect 144362 10996 144368 11008
rect 88300 10968 144368 10996
rect 88300 10956 88306 10968
rect 144362 10956 144368 10968
rect 144420 10956 144426 11008
rect 85666 10276 85672 10328
rect 85724 10316 85730 10328
rect 190638 10316 190644 10328
rect 85724 10288 190644 10316
rect 85724 10276 85730 10288
rect 190638 10276 190644 10288
rect 190696 10276 190702 10328
rect 97902 9596 97908 9648
rect 97960 9636 97966 9648
rect 161566 9636 161572 9648
rect 97960 9608 161572 9636
rect 97960 9596 97966 9608
rect 161566 9596 161572 9608
rect 161624 9596 161630 9648
rect 313274 9596 313280 9648
rect 313332 9636 313338 9648
rect 320818 9636 320824 9648
rect 313332 9608 320824 9636
rect 313332 9596 313338 9608
rect 320818 9596 320824 9608
rect 320876 9596 320882 9648
rect 325602 9596 325608 9648
rect 325660 9636 325666 9648
rect 430666 9636 430672 9648
rect 325660 9608 430672 9636
rect 325660 9596 325666 9608
rect 430666 9596 430672 9608
rect 430724 9596 430730 9648
rect 95142 9528 95148 9580
rect 95200 9568 95206 9580
rect 158438 9568 158444 9580
rect 95200 9540 158444 9568
rect 95200 9528 95206 9540
rect 158438 9528 158444 9540
rect 158496 9528 158502 9580
rect 320726 9528 320732 9580
rect 320784 9568 320790 9580
rect 424410 9568 424416 9580
rect 320784 9540 424416 9568
rect 320784 9528 320790 9540
rect 424410 9528 424416 9540
rect 424468 9528 424474 9580
rect 100754 9460 100760 9512
rect 100812 9500 100818 9512
rect 160002 9500 160008 9512
rect 100812 9472 160008 9500
rect 100812 9460 100818 9472
rect 160002 9460 160008 9472
rect 160060 9460 160066 9512
rect 317322 9460 317328 9512
rect 317380 9500 317386 9512
rect 336182 9500 336188 9512
rect 317380 9472 336188 9500
rect 317380 9460 317386 9472
rect 336182 9460 336188 9472
rect 336240 9460 336246 9512
rect 82814 8236 82820 8288
rect 82872 8276 82878 8288
rect 106826 8276 106832 8288
rect 82872 8248 106832 8276
rect 82872 8236 82878 8248
rect 106826 8236 106832 8248
rect 106884 8236 106890 8288
rect 107654 8236 107660 8288
rect 107712 8276 107718 8288
rect 111518 8276 111524 8288
rect 107712 8248 111524 8276
rect 107712 8236 107718 8248
rect 111518 8236 111524 8248
rect 111576 8236 111582 8288
rect 86862 8168 86868 8220
rect 86920 8208 86926 8220
rect 108390 8208 108396 8220
rect 86920 8180 108396 8208
rect 86920 8168 86926 8180
rect 108390 8168 108396 8180
rect 108448 8168 108454 8220
rect 110414 8168 110420 8220
rect 110472 8208 110478 8220
rect 113082 8208 113088 8220
rect 110472 8180 113088 8208
rect 110472 8168 110478 8180
rect 113082 8168 113088 8180
rect 113140 8168 113146 8220
rect 104802 8100 104808 8152
rect 104860 8140 104866 8152
rect 109954 8140 109960 8152
rect 104860 8112 109960 8140
rect 104860 8100 104866 8112
rect 109954 8100 109960 8112
rect 110012 8100 110018 8152
rect 256694 7828 256700 7880
rect 256752 7868 256758 7880
rect 335538 7868 335544 7880
rect 256752 7840 335544 7868
rect 256752 7828 256758 7840
rect 335538 7828 335544 7840
rect 335596 7828 335602 7880
rect 253198 7692 253204 7744
rect 253256 7732 253262 7744
rect 335722 7732 335728 7744
rect 253256 7704 335728 7732
rect 253256 7692 253262 7704
rect 335722 7692 335728 7704
rect 335780 7692 335786 7744
rect 109310 7624 109316 7676
rect 109368 7664 109374 7676
rect 181898 7664 181904 7676
rect 109368 7636 181904 7664
rect 109368 7624 109374 7636
rect 181898 7624 181904 7636
rect 181956 7624 181962 7676
rect 110506 7556 110512 7608
rect 110564 7596 110570 7608
rect 192110 7596 192116 7608
rect 110564 7568 192116 7596
rect 110564 7556 110570 7568
rect 192110 7556 192116 7568
rect 192168 7556 192174 7608
rect 251082 7556 251088 7608
rect 251140 7596 251146 7608
rect 336090 7596 336096 7608
rect 251140 7568 336096 7596
rect 251140 7556 251146 7568
rect 336090 7556 336096 7568
rect 336148 7556 336154 7608
rect 222102 7352 222108 7404
rect 222160 7392 222166 7404
rect 222838 7392 222844 7404
rect 222160 7364 222844 7392
rect 222160 7352 222166 7364
rect 222838 7352 222844 7364
rect 222896 7352 222902 7404
rect 73154 6808 73160 6860
rect 73212 6848 73218 6860
rect 81802 6848 81808 6860
rect 73212 6820 81808 6848
rect 73212 6808 73218 6820
rect 81802 6808 81808 6820
rect 81860 6808 81866 6860
rect 185670 6808 185676 6860
rect 185728 6848 185734 6860
rect 338574 6848 338580 6860
rect 185728 6820 338580 6848
rect 185728 6808 185734 6820
rect 338574 6808 338580 6820
rect 338632 6808 338638 6860
rect 77202 6740 77208 6792
rect 77260 6780 77266 6792
rect 189810 6780 189816 6792
rect 77260 6752 189816 6780
rect 77260 6740 77266 6752
rect 189810 6740 189816 6752
rect 189868 6740 189874 6792
rect 40678 5448 40684 5500
rect 40736 5488 40742 5500
rect 139670 5488 139676 5500
rect 40736 5460 139676 5488
rect 40736 5448 40742 5460
rect 139670 5448 139676 5460
rect 139728 5448 139734 5500
rect 285582 5448 285588 5500
rect 285640 5488 285646 5500
rect 305638 5488 305644 5500
rect 285640 5460 305644 5488
rect 285640 5448 285646 5460
rect 305638 5448 305644 5460
rect 305696 5448 305702 5500
rect 307662 5448 307668 5500
rect 307720 5488 307726 5500
rect 335906 5488 335912 5500
rect 307720 5460 335912 5488
rect 307720 5448 307726 5460
rect 335906 5448 335912 5460
rect 335964 5448 335970 5500
rect 288434 5380 288440 5432
rect 288492 5420 288498 5432
rect 307018 5420 307024 5432
rect 288492 5392 307024 5420
rect 288492 5380 288498 5392
rect 307018 5380 307024 5392
rect 307076 5380 307082 5432
rect 89714 4836 89720 4888
rect 89772 4876 89778 4888
rect 192662 4876 192668 4888
rect 89772 4848 192668 4876
rect 89772 4836 89778 4848
rect 192662 4836 192668 4848
rect 192720 4836 192726 4888
rect 48958 4768 48964 4820
rect 49016 4808 49022 4820
rect 155310 4808 155316 4820
rect 49016 4780 155316 4808
rect 49016 4768 49022 4780
rect 155310 4768 155316 4780
rect 155368 4768 155374 4820
rect 336642 4768 336648 4820
rect 336700 4808 336706 4820
rect 402514 4808 402520 4820
rect 336700 4780 402520 4808
rect 336700 4768 336706 4780
rect 402514 4768 402520 4780
rect 402572 4768 402578 4820
rect 192110 4196 192116 4208
rect 135180 4168 192116 4196
rect 81434 4088 81440 4140
rect 81492 4128 81498 4140
rect 135180 4128 135208 4168
rect 192110 4156 192116 4168
rect 192168 4156 192174 4208
rect 81492 4100 135208 4128
rect 81492 4088 81498 4100
rect 172422 4088 172428 4140
rect 172480 4128 172486 4140
rect 189902 4128 189908 4140
rect 172480 4100 189908 4128
rect 172480 4088 172486 4100
rect 189902 4088 189908 4100
rect 189960 4088 189966 4140
rect 226426 4088 226432 4140
rect 226484 4128 226490 4140
rect 405642 4128 405648 4140
rect 226484 4100 405648 4128
rect 226484 4088 226490 4100
rect 405642 4088 405648 4100
rect 405700 4088 405706 4140
rect 224954 4020 224960 4072
rect 225012 4060 225018 4072
rect 404078 4060 404084 4072
rect 225012 4032 404084 4060
rect 225012 4020 225018 4032
rect 404078 4020 404084 4032
rect 404136 4020 404142 4072
rect 233878 3952 233884 4004
rect 233936 3992 233942 4004
rect 407206 3992 407212 4004
rect 233936 3964 407212 3992
rect 233936 3952 233942 3964
rect 407206 3952 407212 3964
rect 407264 3952 407270 4004
rect 102134 3544 102140 3596
rect 102192 3584 102198 3596
rect 190822 3584 190828 3596
rect 102192 3556 190828 3584
rect 102192 3544 102198 3556
rect 190822 3544 190828 3556
rect 190880 3544 190886 3596
rect 187326 3476 187332 3528
rect 187384 3516 187390 3528
rect 336642 3516 336648 3528
rect 187384 3488 336648 3516
rect 187384 3476 187390 3488
rect 336642 3476 336648 3488
rect 336700 3476 336706 3528
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 339586 3448 339592 3460
rect 161348 3420 339592 3448
rect 161348 3408 161354 3420
rect 339586 3408 339592 3420
rect 339644 3408 339650 3460
<< via1 >>
rect 338304 85212 338356 85264
rect 338672 85212 338724 85264
rect 337384 80248 337436 80300
rect 336556 80044 336608 80096
rect 336740 80044 336792 80096
rect 337384 80044 337436 80096
rect 81762 79908 81814 79960
rect 398104 79908 398156 79960
rect 338856 79432 338908 79484
rect 338856 79228 338908 79280
rect 124128 78616 124180 78668
rect 173992 78616 174044 78668
rect 178040 78616 178092 78668
rect 329472 78616 329524 78668
rect 118700 78548 118752 78600
rect 152096 78548 152148 78600
rect 117228 78480 117280 78532
rect 142712 78480 142764 78532
rect 320824 78140 320876 78192
rect 400956 78140 401008 78192
rect 305644 78072 305696 78124
rect 408776 78072 408828 78124
rect 174544 78004 174596 78056
rect 302424 78004 302476 78056
rect 307024 78004 307076 78056
rect 411904 78004 411956 78056
rect 181444 77936 181496 77988
rect 333980 77936 334032 77988
rect 144920 77800 144972 77852
rect 146024 77800 146076 77852
rect 75828 12384 75880 12436
rect 191288 12384 191340 12436
rect 78588 12316 78640 12368
rect 191196 12316 191248 12368
rect 88248 10956 88300 11008
rect 144368 10956 144420 11008
rect 85672 10276 85724 10328
rect 190644 10276 190696 10328
rect 97908 9596 97960 9648
rect 161572 9596 161624 9648
rect 313280 9596 313332 9648
rect 320824 9596 320876 9648
rect 325608 9596 325660 9648
rect 430672 9596 430724 9648
rect 95148 9528 95200 9580
rect 158444 9528 158496 9580
rect 320732 9528 320784 9580
rect 424416 9528 424468 9580
rect 100760 9460 100812 9512
rect 160008 9460 160060 9512
rect 317328 9460 317380 9512
rect 336188 9460 336240 9512
rect 82820 8236 82872 8288
rect 106832 8236 106884 8288
rect 107660 8236 107712 8288
rect 111524 8236 111576 8288
rect 86868 8168 86920 8220
rect 108396 8168 108448 8220
rect 110420 8168 110472 8220
rect 113088 8168 113140 8220
rect 104808 8100 104860 8152
rect 109960 8100 110012 8152
rect 256700 7828 256752 7880
rect 335544 7828 335596 7880
rect 253204 7692 253256 7744
rect 335728 7692 335780 7744
rect 109316 7624 109368 7676
rect 181904 7624 181956 7676
rect 110512 7556 110564 7608
rect 192116 7556 192168 7608
rect 251088 7556 251140 7608
rect 336096 7556 336148 7608
rect 222108 7352 222160 7404
rect 222844 7352 222896 7404
rect 73160 6808 73212 6860
rect 81808 6808 81860 6860
rect 185676 6808 185728 6860
rect 338580 6808 338632 6860
rect 77208 6740 77260 6792
rect 189816 6740 189868 6792
rect 40684 5448 40736 5500
rect 139676 5448 139728 5500
rect 285588 5448 285640 5500
rect 305644 5448 305696 5500
rect 307668 5448 307720 5500
rect 335912 5448 335964 5500
rect 288440 5380 288492 5432
rect 307024 5380 307076 5432
rect 89720 4836 89772 4888
rect 192668 4836 192720 4888
rect 48964 4768 49016 4820
rect 155316 4768 155368 4820
rect 336648 4768 336700 4820
rect 402520 4768 402572 4820
rect 81440 4088 81492 4140
rect 192116 4156 192168 4208
rect 172428 4088 172480 4140
rect 189908 4088 189960 4140
rect 226432 4088 226484 4140
rect 405648 4088 405700 4140
rect 224960 4020 225012 4072
rect 404084 4020 404136 4072
rect 233884 3952 233936 4004
rect 407212 3952 407264 4004
rect 102140 3544 102192 3596
rect 190828 3544 190880 3596
rect 187332 3476 187384 3528
rect 336648 3476 336700 3528
rect 161296 3408 161348 3460
rect 339592 3408 339644 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 348804 700505 348832 703520
rect 348790 700496 348846 700505
rect 348790 700431 348846 700440
rect 109038 700360 109094 700369
rect 109038 700295 109094 700304
rect 104714 697232 104770 697241
rect 104714 697167 104770 697176
rect 100390 644056 100446 644065
rect 100390 643991 100446 644000
rect 96066 591016 96122 591025
rect 96066 590951 96122 590960
rect 91742 537840 91798 537849
rect 91742 537775 91798 537784
rect 87418 484664 87474 484673
rect 87418 484599 87474 484608
rect 83094 298752 83150 298761
rect 83094 298687 83150 298696
rect 83108 189938 83136 298687
rect 87432 189938 87460 484599
rect 91756 189938 91784 537775
rect 96080 189938 96108 590951
rect 100404 189938 100432 643991
rect 104728 189938 104756 697167
rect 109052 189938 109080 700295
rect 152278 630864 152334 630873
rect 152278 630799 152334 630808
rect 147954 577688 148010 577697
rect 147954 577623 148010 577632
rect 143630 524512 143686 524521
rect 143630 524447 143686 524456
rect 139306 471472 139362 471481
rect 139306 471407 139362 471416
rect 118054 192672 118110 192681
rect 118054 192607 118110 192616
rect 113638 192536 113694 192545
rect 113638 192471 113694 192480
rect 113652 189938 113680 192471
rect 118068 189938 118096 192607
rect 139320 189938 139348 471407
rect 143644 189938 143672 524447
rect 147968 189938 147996 577623
rect 152292 189938 152320 630799
rect 397472 192681 397500 703520
rect 397458 192672 397514 192681
rect 397458 192607 397514 192616
rect 462332 192545 462360 703520
rect 527192 700369 527220 703520
rect 527178 700360 527234 700369
rect 527178 700295 527234 700304
rect 462318 192536 462374 192545
rect 462318 192471 462374 192480
rect 83076 189910 83136 189938
rect 87400 189910 87460 189938
rect 91724 189910 91784 189938
rect 96048 189910 96108 189938
rect 100372 189910 100432 189938
rect 104696 189910 104756 189938
rect 109020 189910 109080 189938
rect 113344 189910 113680 189938
rect 117668 189910 118096 189938
rect 139288 189910 139348 189938
rect 143612 189910 143672 189938
rect 147936 189910 147996 189938
rect 152260 189910 152320 189938
rect 191838 186552 191894 186561
rect 191838 186487 191894 186496
rect 190458 164656 190514 164665
rect 190458 164591 190514 164600
rect 189998 135824 190054 135833
rect 189998 135759 190054 135768
rect 189354 123448 189410 123457
rect 189354 123383 189410 123392
rect 81774 79966 81802 80036
rect 81762 79960 81814 79966
rect 81762 79902 81814 79908
rect 81774 79778 81802 79902
rect 83338 79778 83366 80036
rect 84902 79778 84930 80036
rect 86466 79778 86494 80036
rect 81774 79750 81848 79778
rect 83338 79750 83412 79778
rect 4066 78024 4122 78033
rect 4066 77959 4122 77968
rect 1674 6624 1730 6633
rect 1674 6559 1730 6568
rect 570 5672 626 5681
rect 570 5607 626 5616
rect 584 480 612 5607
rect 1688 480 1716 6559
rect 2870 3088 2926 3097
rect 2870 3023 2926 3032
rect 2884 480 2912 3023
rect 4080 480 4108 77959
rect 5262 77888 5318 77897
rect 5262 77823 5318 77832
rect 5276 480 5304 77823
rect 41878 77480 41934 77489
rect 41878 77415 41934 77424
rect 18234 77344 18290 77353
rect 18234 77279 18290 77288
rect 7654 6760 7710 6769
rect 7654 6695 7710 6704
rect 6458 3768 6514 3777
rect 6458 3703 6514 3712
rect 6472 480 6500 3703
rect 7668 480 7696 6695
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 9954 5808 10010 5817
rect 9954 5743 10010 5752
rect 8758 4176 8814 4185
rect 8758 4111 8814 4120
rect 8772 480 8800 4111
rect 9968 480 9996 5743
rect 12346 2816 12402 2825
rect 12346 2751 12402 2760
rect 12360 480 12388 2751
rect 13556 480 13584 6151
rect 17038 4856 17094 4865
rect 17038 4791 17094 4800
rect 14738 2952 14794 2961
rect 14738 2887 14794 2896
rect 14752 480 14780 2887
rect 17052 480 17080 4791
rect 18248 480 18276 77279
rect 32402 11112 32458 11121
rect 32402 11047 32458 11056
rect 31298 10296 31354 10305
rect 31298 10231 31354 10240
rect 23018 9752 23074 9761
rect 23018 9687 23074 9696
rect 21822 4992 21878 5001
rect 21822 4927 21878 4936
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19444 480 19472 2751
rect 21836 480 21864 4927
rect 23032 480 23060 9687
rect 30102 5264 30158 5273
rect 30102 5199 30158 5208
rect 26514 5128 26570 5137
rect 26514 5063 26570 5072
rect 24214 3632 24270 3641
rect 24214 3567 24270 3576
rect 24228 480 24256 3567
rect 26528 480 26556 5063
rect 27710 3496 27766 3505
rect 27710 3431 27766 3440
rect 27724 480 27752 3431
rect 28906 3360 28962 3369
rect 28906 3295 28962 3304
rect 28920 480 28948 3295
rect 30116 480 30144 5199
rect 31312 480 31340 10231
rect 32416 480 32444 11047
rect 38382 10568 38438 10577
rect 38382 10503 38438 10512
rect 34794 10432 34850 10441
rect 34794 10367 34850 10376
rect 33598 5400 33654 5409
rect 33598 5335 33654 5344
rect 33612 480 33640 5335
rect 34808 480 34836 10367
rect 37186 5536 37242 5545
rect 37186 5471 37242 5480
rect 35990 3904 36046 3913
rect 35990 3839 36046 3848
rect 36004 480 36032 3839
rect 37200 480 37228 5471
rect 38396 480 38424 10503
rect 40684 5500 40736 5506
rect 40684 5442 40736 5448
rect 40696 4185 40724 5442
rect 40774 4720 40830 4729
rect 40774 4655 40830 4664
rect 40682 4176 40738 4185
rect 40682 4111 40738 4120
rect 40682 4040 40738 4049
rect 40682 3975 40738 3984
rect 40696 3641 40724 3975
rect 40682 3632 40738 3641
rect 40682 3567 40738 3576
rect 39578 3496 39634 3505
rect 39578 3431 39634 3440
rect 39592 480 39620 3431
rect 40788 2394 40816 4655
rect 40696 2366 40816 2394
rect 40696 480 40724 2366
rect 41892 480 41920 77415
rect 67914 13016 67970 13025
rect 67914 12951 67970 12960
rect 64326 12064 64382 12073
rect 64326 11999 64382 12008
rect 60830 11928 60886 11937
rect 60830 11863 60886 11872
rect 53746 11792 53802 11801
rect 53746 11727 53802 11736
rect 50158 11656 50214 11665
rect 50158 11591 50214 11600
rect 46662 11248 46718 11257
rect 46662 11183 46718 11192
rect 45466 10704 45522 10713
rect 45466 10639 45522 10648
rect 44270 9208 44326 9217
rect 44270 9143 44326 9152
rect 43074 3224 43130 3233
rect 43074 3159 43130 3168
rect 43088 480 43116 3159
rect 44284 480 44312 9143
rect 45480 480 45508 10639
rect 46676 480 46704 11183
rect 47858 6896 47914 6905
rect 47858 6831 47914 6840
rect 47872 480 47900 6831
rect 48964 4820 49016 4826
rect 48964 4762 49016 4768
rect 48976 480 49004 4762
rect 50172 480 50200 11591
rect 51354 7440 51410 7449
rect 51354 7375 51410 7384
rect 51368 480 51396 7375
rect 52550 6352 52606 6361
rect 52550 6287 52606 6296
rect 52564 480 52592 6287
rect 53760 480 53788 11727
rect 56046 8528 56102 8537
rect 56046 8463 56102 8472
rect 54942 7984 54998 7993
rect 54942 7919 54998 7928
rect 54956 480 54984 7919
rect 56060 480 56088 8463
rect 59634 8392 59690 8401
rect 59634 8327 59690 8336
rect 58438 7168 58494 7177
rect 58438 7103 58494 7112
rect 57242 3224 57298 3233
rect 57242 3159 57298 3168
rect 57256 480 57284 3159
rect 58452 480 58480 7103
rect 59648 480 59676 8327
rect 60844 480 60872 11863
rect 63222 8664 63278 8673
rect 63222 8599 63278 8608
rect 62026 7032 62082 7041
rect 62026 6967 62082 6976
rect 62040 480 62068 6967
rect 63236 480 63264 8599
rect 64340 480 64368 11999
rect 65522 7304 65578 7313
rect 65522 7239 65578 7248
rect 65536 480 65564 7239
rect 66718 3224 66774 3233
rect 66718 3159 66774 3168
rect 66732 480 66760 3159
rect 67928 480 67956 12951
rect 75828 12436 75880 12442
rect 75828 12378 75880 12384
rect 74998 12336 75054 12345
rect 74998 12271 75054 12280
rect 71502 12200 71558 12209
rect 71502 12135 71558 12144
rect 70306 8936 70362 8945
rect 70306 8871 70362 8880
rect 69110 3224 69166 3233
rect 69110 3159 69166 3168
rect 69124 480 69152 3159
rect 70320 480 70348 8871
rect 71516 480 71544 12135
rect 72606 7576 72662 7585
rect 72606 7511 72662 7520
rect 72620 480 72648 7511
rect 73160 6860 73212 6866
rect 73160 6802 73212 6808
rect 73172 5681 73200 6802
rect 73802 6488 73858 6497
rect 73802 6423 73858 6432
rect 73158 5672 73214 5681
rect 73158 5607 73214 5616
rect 73816 480 73844 6423
rect 75012 480 75040 12271
rect 75840 11121 75868 12378
rect 78588 12368 78640 12374
rect 78588 12310 78640 12316
rect 78494 11520 78550 11529
rect 78494 11455 78550 11464
rect 75826 11112 75882 11121
rect 75826 11047 75882 11056
rect 77390 9072 77446 9081
rect 77390 9007 77446 9016
rect 77208 6792 77260 6798
rect 77208 6734 77260 6740
rect 77220 5817 77248 6734
rect 77206 5808 77262 5817
rect 77206 5743 77262 5752
rect 76194 5672 76250 5681
rect 76194 5607 76250 5616
rect 76208 480 76236 5607
rect 77404 480 77432 9007
rect 78508 6914 78536 11455
rect 78600 11257 78628 12310
rect 78586 11248 78642 11257
rect 78586 11183 78642 11192
rect 80886 10840 80942 10849
rect 80886 10775 80942 10784
rect 79690 7712 79746 7721
rect 79690 7647 79746 7656
rect 78508 6886 78628 6914
rect 78600 480 78628 6886
rect 79704 480 79732 7647
rect 80900 480 80928 10775
rect 81820 6866 81848 79750
rect 82820 8288 82872 8294
rect 82820 8230 82872 8236
rect 82832 7449 82860 8230
rect 83094 7848 83150 7857
rect 83094 7783 83150 7792
rect 83278 7848 83334 7857
rect 83278 7783 83334 7792
rect 83108 7449 83136 7783
rect 82818 7440 82874 7449
rect 82818 7375 82874 7384
rect 83094 7440 83150 7449
rect 83094 7375 83150 7384
rect 81808 6860 81860 6866
rect 81808 6802 81860 6808
rect 81440 4140 81492 4146
rect 81440 4082 81492 4088
rect 81452 3097 81480 4082
rect 82082 3224 82138 3233
rect 82082 3159 82138 3168
rect 81438 3088 81494 3097
rect 81438 3023 81494 3032
rect 82096 480 82124 3159
rect 83292 480 83320 7783
rect 83384 6633 83412 79750
rect 84856 79750 84930 79778
rect 86420 79750 86494 79778
rect 88030 79778 88058 80036
rect 89594 79778 89622 80036
rect 91158 79778 91186 80036
rect 88030 79750 88104 79778
rect 89594 79750 89668 79778
rect 84856 78033 84884 79750
rect 84842 78024 84898 78033
rect 84842 77959 84898 77968
rect 86420 77897 86448 79750
rect 86406 77888 86462 77897
rect 86406 77823 86462 77832
rect 84474 10976 84530 10985
rect 84474 10911 84530 10920
rect 83370 6624 83426 6633
rect 83370 6559 83426 6568
rect 84488 480 84516 10911
rect 85672 10328 85724 10334
rect 85672 10270 85724 10276
rect 85684 480 85712 10270
rect 87970 10160 88026 10169
rect 87970 10095 88026 10104
rect 86868 8220 86920 8226
rect 86868 8162 86920 8168
rect 86880 7993 86908 8162
rect 86866 7984 86922 7993
rect 87050 7984 87106 7993
rect 86866 7919 86922 7928
rect 86972 7942 87050 7970
rect 86972 7834 87000 7942
rect 87050 7919 87106 7928
rect 86880 7806 87000 7834
rect 86880 480 86908 7806
rect 87984 480 88012 10095
rect 88076 3641 88104 79750
rect 88248 11008 88300 11014
rect 88248 10950 88300 10956
rect 88260 9761 88288 10950
rect 88246 9752 88302 9761
rect 88246 9687 88302 9696
rect 89640 6769 89668 79750
rect 91112 79750 91186 79778
rect 92722 79778 92750 80036
rect 94286 79778 94314 80036
rect 95850 79778 95878 80036
rect 97414 79778 97442 80036
rect 98978 79778 99006 80036
rect 100542 79778 100570 80036
rect 102106 79778 102134 80036
rect 103670 79778 103698 80036
rect 105234 79778 105262 80036
rect 106798 79778 106826 80036
rect 108362 79778 108390 80036
rect 109926 79778 109954 80036
rect 111490 79778 111518 80036
rect 113054 79778 113082 80036
rect 114618 79778 114646 80036
rect 116182 79778 116210 80036
rect 117746 79778 117774 80036
rect 119310 79778 119338 80036
rect 120874 79778 120902 80036
rect 122438 79778 122466 80036
rect 124002 79778 124030 80036
rect 125566 79778 125594 80036
rect 127130 79778 127158 80036
rect 128694 79778 128722 80036
rect 130258 79778 130286 80036
rect 131822 79778 131850 80036
rect 133386 79778 133414 80036
rect 134950 79778 134978 80036
rect 136514 79778 136542 80036
rect 138078 79778 138106 80036
rect 139642 79778 139670 80036
rect 141206 79778 141234 80036
rect 142770 79778 142798 80036
rect 92722 79750 92796 79778
rect 94286 79750 94360 79778
rect 95850 79750 95924 79778
rect 97414 79750 97488 79778
rect 98978 79750 99052 79778
rect 100542 79750 100616 79778
rect 102106 79750 102180 79778
rect 103670 79750 103744 79778
rect 105234 79750 105308 79778
rect 106798 79750 106872 79778
rect 108362 79750 108436 79778
rect 109926 79750 110000 79778
rect 111490 79750 111564 79778
rect 113054 79750 113128 79778
rect 114618 79750 114692 79778
rect 116182 79750 116256 79778
rect 117746 79750 117820 79778
rect 119310 79750 119384 79778
rect 120874 79750 120948 79778
rect 122438 79750 122512 79778
rect 124002 79750 124076 79778
rect 125566 79750 125640 79778
rect 127130 79750 127204 79778
rect 128694 79750 128768 79778
rect 130258 79750 130332 79778
rect 131822 79750 131896 79778
rect 133386 79750 133460 79778
rect 134950 79750 135024 79778
rect 136514 79750 136588 79778
rect 138078 79750 138152 79778
rect 139642 79750 139716 79778
rect 141206 79750 141280 79778
rect 91112 77353 91140 79750
rect 91558 78296 91614 78305
rect 91558 78231 91614 78240
rect 91098 77344 91154 77353
rect 91098 77279 91154 77288
rect 90362 9344 90418 9353
rect 90362 9279 90418 9288
rect 89626 6760 89682 6769
rect 89626 6695 89682 6704
rect 89166 6624 89222 6633
rect 89166 6559 89222 6568
rect 88062 3632 88118 3641
rect 88062 3567 88118 3576
rect 88982 3632 89038 3641
rect 88982 3567 89038 3576
rect 88996 3233 89024 3567
rect 88982 3224 89038 3233
rect 88982 3159 89038 3168
rect 89180 480 89208 6559
rect 89720 4888 89772 4894
rect 89720 4830 89772 4836
rect 89732 3913 89760 4830
rect 89718 3904 89774 3913
rect 89718 3839 89774 3848
rect 90376 480 90404 9279
rect 91572 480 91600 78231
rect 92768 6914 92796 79750
rect 93950 9480 94006 9489
rect 93950 9415 94006 9424
rect 92676 6886 92796 6914
rect 92676 4865 92704 6886
rect 92754 6760 92810 6769
rect 92754 6695 92810 6704
rect 92662 4856 92718 4865
rect 92662 4791 92718 4800
rect 92768 480 92796 6695
rect 93964 480 93992 9415
rect 94332 5001 94360 79750
rect 95148 9580 95200 9586
rect 95148 9522 95200 9528
rect 95160 8537 95188 9522
rect 95146 8528 95202 8537
rect 95146 8463 95202 8472
rect 95896 5137 95924 79750
rect 97460 5273 97488 79750
rect 98642 77888 98698 77897
rect 98642 77823 98698 77832
rect 98656 16574 98684 77823
rect 98472 16546 98684 16574
rect 97908 9648 97960 9654
rect 97814 9616 97870 9625
rect 97908 9590 97960 9596
rect 97814 9551 97870 9560
rect 97446 5264 97502 5273
rect 97446 5199 97502 5208
rect 95882 5128 95938 5137
rect 95882 5063 95938 5072
rect 94318 4992 94374 5001
rect 94318 4927 94374 4936
rect 95146 3768 95202 3777
rect 95146 3703 95202 3712
rect 96250 3768 96306 3777
rect 96250 3703 96306 3712
rect 95160 480 95188 3703
rect 96264 480 96292 3703
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 354 97530 480
rect 97828 354 97856 9551
rect 97920 8673 97948 9590
rect 97906 8664 97962 8673
rect 97906 8599 97962 8608
rect 98472 6914 98500 16546
rect 98550 7440 98606 7449
rect 98550 7375 98606 7384
rect 98564 7154 98592 7375
rect 98826 7168 98882 7177
rect 98564 7126 98826 7154
rect 98826 7103 98882 7112
rect 98472 6886 98684 6914
rect 98656 480 98684 6886
rect 99024 5409 99052 79750
rect 100588 5545 100616 79750
rect 100760 9512 100812 9518
rect 100760 9454 100812 9460
rect 100772 8401 100800 9454
rect 101034 8800 101090 8809
rect 101034 8735 101090 8744
rect 100758 8392 100814 8401
rect 100758 8327 100814 8336
rect 100574 5536 100630 5545
rect 100574 5471 100630 5480
rect 99010 5400 99066 5409
rect 99010 5335 99066 5344
rect 99838 4040 99894 4049
rect 99838 3975 99894 3984
rect 99852 480 99880 3975
rect 101048 480 101076 8735
rect 102152 4729 102180 79750
rect 102230 78024 102286 78033
rect 102230 77959 102286 77968
rect 102138 4720 102194 4729
rect 102138 4655 102194 4664
rect 102140 3596 102192 3602
rect 102140 3538 102192 3544
rect 102152 2961 102180 3538
rect 102138 2952 102194 2961
rect 102138 2887 102194 2896
rect 102244 480 102272 77959
rect 103716 9217 103744 79750
rect 103702 9208 103758 9217
rect 103702 9143 103758 9152
rect 104808 8152 104860 8158
rect 104530 8120 104586 8129
rect 104808 8094 104860 8100
rect 104530 8055 104586 8064
rect 103334 3224 103390 3233
rect 103334 3159 103390 3168
rect 103348 480 103376 3159
rect 104544 480 104572 8055
rect 104820 7449 104848 8094
rect 104806 7440 104862 7449
rect 104806 7375 104862 7384
rect 105280 6905 105308 79750
rect 105726 78568 105782 78577
rect 105726 78503 105782 78512
rect 105266 6896 105322 6905
rect 105266 6831 105322 6840
rect 105740 480 105768 78503
rect 106844 8294 106872 79750
rect 106832 8288 106884 8294
rect 106832 8230 106884 8236
rect 107660 8288 107712 8294
rect 107660 8230 107712 8236
rect 108118 8256 108174 8265
rect 107672 7041 107700 8230
rect 108408 8226 108436 79750
rect 108118 8191 108174 8200
rect 108396 8220 108448 8226
rect 107658 7032 107714 7041
rect 107658 6967 107714 6976
rect 106922 6896 106978 6905
rect 106922 6831 106978 6840
rect 106936 480 106964 6831
rect 108132 480 108160 8191
rect 108396 8162 108448 8168
rect 109972 8158 110000 79750
rect 111536 8294 111564 79750
rect 112810 77752 112866 77761
rect 112810 77687 112866 77696
rect 111524 8288 111576 8294
rect 111524 8230 111576 8236
rect 110420 8220 110472 8226
rect 110420 8162 110472 8168
rect 109960 8152 110012 8158
rect 109960 8094 110012 8100
rect 109316 7676 109368 7682
rect 109316 7618 109368 7624
rect 109328 480 109356 7618
rect 110432 7313 110460 8162
rect 110512 7608 110564 7614
rect 110512 7550 110564 7556
rect 110418 7304 110474 7313
rect 110418 7239 110474 7248
rect 110524 480 110552 7550
rect 111614 7440 111670 7449
rect 111614 7375 111670 7384
rect 111628 480 111656 7375
rect 112824 480 112852 77687
rect 113100 8226 113128 79750
rect 114664 77353 114692 79750
rect 116122 78160 116178 78169
rect 116122 78095 116178 78104
rect 116136 77625 116164 78095
rect 116122 77616 116178 77625
rect 116122 77551 116178 77560
rect 114650 77344 114706 77353
rect 114650 77279 114706 77288
rect 113088 8220 113140 8226
rect 113088 8162 113140 8168
rect 116228 7585 116256 79750
rect 117228 78532 117280 78538
rect 117228 78474 117280 78480
rect 116398 77616 116454 77625
rect 116398 77551 116454 77560
rect 116214 7576 116270 7585
rect 116214 7511 116270 7520
rect 115202 4856 115258 4865
rect 115202 4791 115258 4800
rect 114006 2952 114062 2961
rect 114006 2887 114062 2896
rect 114020 480 114048 2887
rect 115216 480 115244 4791
rect 116412 480 116440 77551
rect 117240 77489 117268 78474
rect 117226 77480 117282 77489
rect 117226 77415 117282 77424
rect 117792 6089 117820 79750
rect 118700 78600 118752 78606
rect 118700 78542 118752 78548
rect 118712 78169 118740 78542
rect 118698 78160 118754 78169
rect 118698 78095 118754 78104
rect 119356 7721 119384 79750
rect 119894 77480 119950 77489
rect 119894 77415 119950 77424
rect 119342 7712 119398 7721
rect 119342 7647 119398 7656
rect 117778 6080 117834 6089
rect 117778 6015 117834 6024
rect 118790 5400 118846 5409
rect 118790 5335 118846 5344
rect 117594 4992 117650 5001
rect 117594 4927 117650 4936
rect 117608 480 117636 4927
rect 118804 480 118832 5335
rect 119908 480 119936 77415
rect 120920 7857 120948 79750
rect 122484 7993 122512 79750
rect 123482 77344 123538 77353
rect 123482 77279 123538 77288
rect 122470 7984 122526 7993
rect 122470 7919 122526 7928
rect 120906 7848 120962 7857
rect 120906 7783 120962 7792
rect 122286 5536 122342 5545
rect 122286 5471 122342 5480
rect 121090 5128 121146 5137
rect 121090 5063 121146 5072
rect 121104 480 121132 5063
rect 122300 480 122328 5471
rect 123496 480 123524 77279
rect 124048 9353 124076 79750
rect 124128 78668 124180 78674
rect 124128 78610 124180 78616
rect 124140 78305 124168 78610
rect 124126 78296 124182 78305
rect 124126 78231 124182 78240
rect 125612 9489 125640 79750
rect 127176 9625 127204 79750
rect 127162 9616 127218 9625
rect 127162 9551 127218 9560
rect 125598 9480 125654 9489
rect 125598 9415 125654 9424
rect 124034 9344 124090 9353
rect 124034 9279 124090 9288
rect 128740 8809 128768 79750
rect 128726 8800 128782 8809
rect 128726 8735 128782 8744
rect 130304 8129 130332 79750
rect 131868 8265 131896 79750
rect 131854 8256 131910 8265
rect 131854 8191 131910 8200
rect 130290 8120 130346 8129
rect 130290 8055 130346 8064
rect 133432 7449 133460 79750
rect 133418 7440 133474 7449
rect 133418 7375 133474 7384
rect 124678 5264 124734 5273
rect 124678 5199 124734 5208
rect 124692 480 124720 5199
rect 134996 4865 135024 79750
rect 136560 5409 136588 79750
rect 138124 5545 138152 79750
rect 138110 5536 138166 5545
rect 139688 5506 139716 79750
rect 141252 6225 141280 79750
rect 142724 79750 142798 79778
rect 144334 79778 144362 80036
rect 145898 79778 145926 80036
rect 144334 79750 144408 79778
rect 142724 78538 142752 79750
rect 142712 78532 142764 78538
rect 142712 78474 142764 78480
rect 144380 11014 144408 79750
rect 145852 79750 145926 79778
rect 147462 79778 147490 80036
rect 149026 79778 149054 80036
rect 150590 79778 150618 80036
rect 152154 79778 152182 80036
rect 147462 79750 147536 79778
rect 149026 79750 149100 79778
rect 150590 79750 150664 79778
rect 145852 77897 145880 79750
rect 144918 77888 144974 77897
rect 144918 77823 144920 77832
rect 144972 77823 144974 77832
rect 145838 77888 145894 77897
rect 145838 77823 145894 77832
rect 146022 77888 146078 77897
rect 146022 77823 146024 77832
rect 144920 77794 144972 77800
rect 146076 77823 146078 77832
rect 146024 77794 146076 77800
rect 144368 11008 144420 11014
rect 144368 10950 144420 10956
rect 147508 10305 147536 79750
rect 149072 10441 149100 79750
rect 150636 10577 150664 79750
rect 152108 79750 152182 79778
rect 153718 79778 153746 80036
rect 155282 79778 155310 80036
rect 156846 79778 156874 80036
rect 158410 79778 158438 80036
rect 159974 79778 160002 80036
rect 161538 79778 161566 80036
rect 163102 79778 163130 80036
rect 153718 79750 153792 79778
rect 155282 79750 155356 79778
rect 156846 79750 156920 79778
rect 158410 79750 158484 79778
rect 159974 79750 160048 79778
rect 161538 79750 161612 79778
rect 152108 78606 152136 79750
rect 152096 78600 152148 78606
rect 152096 78542 152148 78548
rect 153764 10713 153792 79750
rect 153750 10704 153806 10713
rect 153750 10639 153806 10648
rect 150622 10568 150678 10577
rect 150622 10503 150678 10512
rect 149058 10432 149114 10441
rect 149058 10367 149114 10376
rect 147494 10296 147550 10305
rect 147494 10231 147550 10240
rect 154210 7712 154266 7721
rect 154210 7647 154266 7656
rect 141238 6216 141294 6225
rect 141238 6151 141294 6160
rect 138110 5471 138166 5480
rect 139676 5500 139728 5506
rect 139676 5442 139728 5448
rect 136546 5400 136602 5409
rect 136546 5335 136602 5344
rect 134982 4856 135038 4865
rect 134982 4791 135038 4800
rect 154224 480 154252 7647
rect 155328 4826 155356 79750
rect 155406 8392 155462 8401
rect 155406 8327 155462 8336
rect 155316 4820 155368 4826
rect 155316 4762 155368 4768
rect 155420 480 155448 8327
rect 156892 6361 156920 79750
rect 158456 9586 158484 79750
rect 158902 10296 158958 10305
rect 158902 10231 158958 10240
rect 158444 9580 158496 9586
rect 158444 9522 158496 9528
rect 156878 6352 156934 6361
rect 156878 6287 156934 6296
rect 157798 5672 157854 5681
rect 157798 5607 157854 5616
rect 156602 5400 156658 5409
rect 156602 5335 156658 5344
rect 156616 480 156644 5335
rect 157812 480 157840 5607
rect 158916 480 158944 10231
rect 160020 9518 160048 79750
rect 161584 9654 161612 79750
rect 163056 79750 163130 79778
rect 164666 79778 164694 80036
rect 166230 79778 166258 80036
rect 167794 79778 167822 80036
rect 169358 79778 169386 80036
rect 170922 79778 170950 80036
rect 172486 79778 172514 80036
rect 174050 79778 174078 80036
rect 175614 79778 175642 80036
rect 177178 79778 177206 80036
rect 178742 79778 178770 80036
rect 180306 79778 180334 80036
rect 164666 79750 164740 79778
rect 166230 79750 166304 79778
rect 167794 79750 167868 79778
rect 169358 79750 169432 79778
rect 170922 79750 170996 79778
rect 172486 79750 172560 79778
rect 163056 78169 163084 79750
rect 163042 78160 163098 78169
rect 163042 78095 163098 78104
rect 161572 9648 161624 9654
rect 161572 9590 161624 9596
rect 160008 9512 160060 9518
rect 160008 9454 160060 9460
rect 164712 8945 164740 79750
rect 164882 10432 164938 10441
rect 164882 10367 164938 10376
rect 164698 8936 164754 8945
rect 164698 8871 164754 8880
rect 162490 7032 162546 7041
rect 162490 6967 162546 6976
rect 160098 6352 160154 6361
rect 160098 6287 160154 6296
rect 160112 480 160140 6287
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 161308 480 161336 3402
rect 162504 480 162532 6967
rect 163686 4856 163742 4865
rect 163686 4791 163742 4800
rect 163700 480 163728 4791
rect 164896 480 164924 10367
rect 166078 7168 166134 7177
rect 166078 7103 166134 7112
rect 166092 480 166120 7103
rect 166276 6497 166304 79750
rect 167840 9081 167868 79750
rect 168378 79384 168434 79393
rect 168378 79319 168434 79328
rect 167826 9072 167882 9081
rect 167826 9007 167882 9016
rect 166262 6488 166318 6497
rect 166262 6423 166318 6432
rect 167182 5536 167238 5545
rect 167182 5471 167238 5480
rect 167196 480 167224 5471
rect 168392 480 168420 79319
rect 169404 10849 169432 79750
rect 170968 10985 170996 79750
rect 170954 10976 171010 10985
rect 170954 10911 171010 10920
rect 169390 10840 169446 10849
rect 169390 10775 169446 10784
rect 172532 10169 172560 79750
rect 174004 79750 174078 79778
rect 175568 79750 175642 79778
rect 177132 79750 177206 79778
rect 178696 79750 178770 79778
rect 180260 79750 180334 79778
rect 181870 79778 181898 80036
rect 183434 79778 183462 80036
rect 184998 79778 185026 80036
rect 186562 79778 186590 80036
rect 188126 79778 188154 80036
rect 181870 79750 181944 79778
rect 174004 78674 174032 79750
rect 173992 78668 174044 78674
rect 173992 78610 174044 78616
rect 174544 78056 174596 78062
rect 174544 77998 174596 78004
rect 172518 10160 172574 10169
rect 172518 10095 172574 10104
rect 169574 7576 169630 7585
rect 169574 7511 169630 7520
rect 169588 480 169616 7511
rect 174556 5409 174584 77998
rect 175568 77897 175596 79750
rect 177132 78033 177160 79750
rect 178040 78668 178092 78674
rect 178040 78610 178092 78616
rect 177118 78024 177174 78033
rect 177118 77959 177174 77968
rect 175554 77888 175610 77897
rect 175554 77823 175610 77832
rect 178052 77330 178080 78610
rect 178696 78441 178724 79750
rect 180260 78577 180288 79750
rect 180246 78568 180302 78577
rect 180246 78503 180302 78512
rect 178682 78432 178738 78441
rect 178682 78367 178738 78376
rect 179234 78432 179290 78441
rect 179234 78367 179290 78376
rect 178958 78160 179014 78169
rect 178958 78095 179014 78104
rect 177868 77302 178080 77330
rect 175462 6216 175518 6225
rect 175462 6151 175518 6160
rect 174542 5400 174598 5409
rect 174542 5335 174598 5344
rect 170770 4720 170826 4729
rect 170770 4655 170826 4664
rect 170784 480 170812 4655
rect 172978 4312 173034 4321
rect 172978 4247 173034 4256
rect 172428 4140 172480 4146
rect 172428 4082 172480 4088
rect 171966 3088 172022 3097
rect 171966 3023 172022 3032
rect 171980 480 172008 3023
rect 172440 2825 172468 4082
rect 172992 3913 173020 4247
rect 174266 4176 174322 4185
rect 174266 4111 174322 4120
rect 172978 3904 173034 3913
rect 172978 3839 173034 3848
rect 173162 3904 173218 3913
rect 173162 3839 173218 3848
rect 173622 3904 173678 3913
rect 173622 3839 173678 3848
rect 172426 2816 172482 2825
rect 172426 2751 172482 2760
rect 173176 480 173204 3839
rect 173636 3097 173664 3839
rect 173622 3088 173678 3097
rect 173622 3023 173678 3032
rect 174280 480 174308 4111
rect 175476 480 175504 6151
rect 176658 4448 176714 4457
rect 176658 4383 176714 4392
rect 176672 480 176700 4383
rect 177868 480 177896 77302
rect 178972 4729 179000 78095
rect 179248 6361 179276 78367
rect 180062 78296 180118 78305
rect 180062 78231 180118 78240
rect 179234 6352 179290 6361
rect 179234 6287 179290 6296
rect 179050 5808 179106 5817
rect 179050 5743 179106 5752
rect 178958 4720 179014 4729
rect 178958 4655 179014 4664
rect 179064 480 179092 5743
rect 180076 5545 180104 78231
rect 181444 77988 181496 77994
rect 181444 77930 181496 77936
rect 180246 7440 180302 7449
rect 181074 7440 181130 7449
rect 180246 7375 180302 7384
rect 180812 7398 181074 7426
rect 180062 5536 180118 5545
rect 180062 5471 180118 5480
rect 180260 480 180288 7375
rect 180812 7313 180840 7398
rect 181074 7375 181130 7384
rect 180798 7304 180854 7313
rect 180798 7239 180854 7248
rect 181456 480 181484 77930
rect 181916 7682 181944 79750
rect 183388 79750 183462 79778
rect 184952 79750 185026 79778
rect 186516 79750 186590 79778
rect 188080 79750 188154 79778
rect 183388 77761 183416 79750
rect 183374 77752 183430 77761
rect 183374 77687 183430 77696
rect 184952 77625 184980 79750
rect 184938 77616 184994 77625
rect 184938 77551 184994 77560
rect 186516 77489 186544 79750
rect 186502 77480 186558 77489
rect 186502 77415 186558 77424
rect 188080 77353 188108 79750
rect 188066 77344 188122 77353
rect 188066 77279 188122 77288
rect 189368 11801 189396 123383
rect 189446 120320 189502 120329
rect 189446 120255 189502 120264
rect 189354 11792 189410 11801
rect 189354 11727 189410 11736
rect 189460 11665 189488 120255
rect 189538 110936 189594 110945
rect 189538 110871 189594 110880
rect 189446 11656 189502 11665
rect 189446 11591 189502 11600
rect 183742 8528 183798 8537
rect 183742 8463 183798 8472
rect 181904 7676 181956 7682
rect 181904 7618 181956 7624
rect 182546 6352 182602 6361
rect 182546 6287 182602 6296
rect 182560 480 182588 6287
rect 183756 480 183784 8463
rect 185676 6860 185728 6866
rect 185676 6802 185728 6808
rect 185582 6488 185638 6497
rect 185582 6423 185638 6432
rect 185596 6089 185624 6423
rect 185582 6080 185638 6089
rect 185582 6015 185638 6024
rect 185688 5681 185716 6802
rect 186134 6488 186190 6497
rect 186134 6423 186190 6432
rect 185674 5672 185730 5681
rect 185674 5607 185730 5616
rect 185582 3496 185638 3505
rect 185582 3431 185638 3440
rect 185030 3360 185086 3369
rect 185030 3295 185086 3304
rect 185044 2961 185072 3295
rect 185596 3097 185624 3431
rect 185582 3088 185638 3097
rect 185582 3023 185638 3032
rect 185030 2952 185086 2961
rect 185030 2887 185086 2896
rect 186148 480 186176 6423
rect 187332 3528 187384 3534
rect 189552 3505 189580 110871
rect 189630 101552 189686 101561
rect 189630 101487 189686 101496
rect 187332 3470 187384 3476
rect 189538 3496 189594 3505
rect 187344 480 187372 3470
rect 189538 3431 189594 3440
rect 189644 2961 189672 101487
rect 189906 95296 189962 95305
rect 189906 95231 189962 95240
rect 189814 88904 189870 88913
rect 189814 88839 189870 88848
rect 189722 80608 189778 80617
rect 189722 80543 189778 80552
rect 189736 7721 189764 80543
rect 189722 7712 189778 7721
rect 189722 7647 189778 7656
rect 189828 6798 189856 88839
rect 189816 6792 189868 6798
rect 189816 6734 189868 6740
rect 189920 4146 189948 95231
rect 190012 13025 190040 135759
rect 189998 13016 190054 13025
rect 189998 12951 190054 12960
rect 189908 4140 189960 4146
rect 189908 4082 189960 4088
rect 190472 4049 190500 164591
rect 190550 161528 190606 161537
rect 190550 161463 190606 161472
rect 190458 4040 190514 4049
rect 190458 3975 190514 3984
rect 190564 3777 190592 161463
rect 190642 152144 190698 152153
rect 190642 152079 190698 152088
rect 190656 10334 190684 152079
rect 190734 145888 190790 145897
rect 190734 145823 190790 145832
rect 190748 11529 190776 145823
rect 190826 142760 190882 142769
rect 190826 142695 190882 142704
rect 190840 12345 190868 142695
rect 190918 139632 190974 139641
rect 190918 139567 190974 139576
rect 190826 12336 190882 12345
rect 190826 12271 190882 12280
rect 190932 12209 190960 139567
rect 191010 133376 191066 133385
rect 191010 133311 191066 133320
rect 190918 12200 190974 12209
rect 190918 12135 190974 12144
rect 191024 12073 191052 133311
rect 191102 130248 191158 130257
rect 191102 130183 191158 130192
rect 191010 12064 191066 12073
rect 191010 11999 191066 12008
rect 191116 11937 191144 130183
rect 191194 117736 191250 117745
rect 191194 117671 191250 117680
rect 191208 12374 191236 117671
rect 191286 105224 191342 105233
rect 191286 105159 191342 105168
rect 191300 12442 191328 105159
rect 191288 12436 191340 12442
rect 191288 12378 191340 12384
rect 191196 12368 191248 12374
rect 191196 12310 191248 12316
rect 191102 11928 191158 11937
rect 191102 11863 191158 11872
rect 190734 11520 190790 11529
rect 190734 11455 190790 11464
rect 190644 10328 190696 10334
rect 190644 10270 190696 10276
rect 191852 5273 191880 186487
rect 191930 183424 191986 183433
rect 191930 183359 191986 183368
rect 191838 5264 191894 5273
rect 191838 5199 191894 5208
rect 191944 5137 191972 183359
rect 192022 180296 192078 180305
rect 192022 180231 192078 180240
rect 191930 5128 191986 5137
rect 191930 5063 191986 5072
rect 192036 5001 192064 180231
rect 192114 174040 192170 174049
rect 192114 173975 192170 173984
rect 192128 7614 192156 173975
rect 192206 170912 192262 170921
rect 192206 170847 192262 170856
rect 192116 7608 192168 7614
rect 192116 7550 192168 7556
rect 192220 6905 192248 170847
rect 192298 167784 192354 167793
rect 192298 167719 192354 167728
rect 192206 6896 192262 6905
rect 192206 6831 192262 6840
rect 192114 5536 192170 5545
rect 192114 5471 192170 5480
rect 192022 4992 192078 5001
rect 192022 4927 192078 4936
rect 192128 4214 192156 5471
rect 192116 4208 192168 4214
rect 192116 4150 192168 4156
rect 190826 4040 190882 4049
rect 190826 3975 190882 3984
rect 190550 3768 190606 3777
rect 190550 3703 190606 3712
rect 190840 3602 190868 3975
rect 190828 3596 190880 3602
rect 190828 3538 190880 3544
rect 189722 3496 189778 3505
rect 189722 3431 189778 3440
rect 189630 2952 189686 2961
rect 189630 2887 189686 2896
rect 189736 480 189764 3431
rect 192312 3233 192340 167719
rect 192390 158400 192446 158409
rect 192390 158335 192446 158344
rect 192404 6633 192432 158335
rect 192482 155272 192538 155281
rect 192482 155207 192538 155216
rect 192390 6624 192446 6633
rect 192390 6559 192446 6568
rect 192496 6089 192524 155207
rect 192574 149016 192630 149025
rect 192574 148951 192630 148960
rect 192482 6080 192538 6089
rect 192482 6015 192538 6024
rect 192298 3224 192354 3233
rect 192298 3159 192354 3168
rect 192588 3097 192616 148951
rect 267738 120592 267794 120601
rect 267738 120527 267794 120536
rect 304538 120592 304594 120601
rect 304538 120527 304594 120536
rect 264150 120184 264206 120193
rect 264150 120119 264206 120128
rect 192666 108352 192722 108361
rect 192666 108287 192722 108296
rect 192680 4894 192708 108287
rect 193862 80744 193918 80753
rect 193862 80679 193918 80688
rect 192668 4888 192720 4894
rect 192668 4830 192720 4836
rect 193218 4040 193274 4049
rect 193218 3975 193274 3984
rect 192574 3088 192630 3097
rect 192574 3023 192630 3032
rect 190826 2952 190882 2961
rect 190826 2887 190882 2896
rect 190840 480 190868 2887
rect 193232 480 193260 3975
rect 193876 3505 193904 80679
rect 246394 79656 246450 79665
rect 246394 79591 246450 79600
rect 207386 79520 207442 79529
rect 207386 79455 207442 79464
rect 200302 5536 200358 5545
rect 200302 5471 200358 5480
rect 196806 5264 196862 5273
rect 196806 5199 196862 5208
rect 193862 3496 193918 3505
rect 193862 3431 193918 3440
rect 194414 3088 194470 3097
rect 194414 3023 194470 3032
rect 194428 480 194456 3023
rect 196820 480 196848 5199
rect 197910 2816 197966 2825
rect 197910 2751 197966 2760
rect 197924 480 197952 2751
rect 200316 480 200344 5471
rect 201498 4312 201554 4321
rect 201498 4247 201554 4256
rect 201512 480 201540 4247
rect 205086 3768 205142 3777
rect 205086 3703 205142 3712
rect 203890 3224 203946 3233
rect 203890 3159 203946 3168
rect 203904 480 203932 3159
rect 205100 480 205128 3703
rect 207400 480 207428 79455
rect 222750 78024 222806 78033
rect 222750 77959 222806 77968
rect 215666 77888 215722 77897
rect 215666 77823 215722 77832
rect 210974 77616 211030 77625
rect 210974 77551 211030 77560
rect 208582 4448 208638 4457
rect 208582 4383 208638 4392
rect 208596 480 208624 4383
rect 210988 480 211016 77551
rect 214470 6624 214526 6633
rect 214470 6559 214526 6568
rect 212170 3360 212226 3369
rect 212170 3295 212226 3304
rect 212184 480 212212 3295
rect 214484 480 214512 6559
rect 215680 480 215708 77823
rect 218058 22672 218114 22681
rect 218058 22607 218114 22616
rect 218072 480 218100 22607
rect 222108 7404 222160 7410
rect 222108 7346 222160 7352
rect 222120 7041 222148 7346
rect 222106 7032 222162 7041
rect 222106 6967 222162 6976
rect 221554 6760 221610 6769
rect 221554 6695 221610 6704
rect 219254 3632 219310 3641
rect 219254 3567 219310 3576
rect 219268 480 219296 3567
rect 221568 480 221596 6695
rect 222764 480 222792 77959
rect 229834 9072 229890 9081
rect 229834 9007 229890 9016
rect 222842 7440 222898 7449
rect 222842 7375 222844 7384
rect 222896 7375 222898 7384
rect 222844 7346 222896 7352
rect 228730 6896 228786 6905
rect 228730 6831 228786 6840
rect 226432 4140 226484 4146
rect 226432 4082 226484 4088
rect 224960 4072 225012 4078
rect 224960 4014 225012 4020
rect 224972 2961 225000 4014
rect 226338 3496 226394 3505
rect 226338 3431 226394 3440
rect 225142 3224 225198 3233
rect 225142 3159 225198 3168
rect 224958 2952 225014 2961
rect 224958 2887 225014 2896
rect 225156 480 225184 3159
rect 226352 480 226380 3431
rect 226444 3097 226472 4082
rect 226430 3088 226486 3097
rect 226430 3023 226486 3032
rect 228744 480 228772 6831
rect 229848 480 229876 9007
rect 242898 7984 242954 7993
rect 242898 7919 242954 7928
rect 239310 7848 239366 7857
rect 239310 7783 239366 7792
rect 235814 7712 235870 7721
rect 235814 7647 235870 7656
rect 232226 6080 232282 6089
rect 232226 6015 232282 6024
rect 232240 480 232268 6015
rect 233884 4004 233936 4010
rect 233884 3946 233936 3952
rect 233238 3768 233294 3777
rect 233238 3703 233294 3712
rect 233422 3768 233478 3777
rect 233422 3703 233478 3712
rect 233252 2961 233280 3703
rect 233238 2952 233294 2961
rect 233238 2887 233294 2896
rect 233436 480 233464 3703
rect 233896 2825 233924 3946
rect 233882 2816 233938 2825
rect 233882 2751 233938 2760
rect 235828 480 235856 7647
rect 239324 480 239352 7783
rect 242912 480 242940 7919
rect 243358 7440 243414 7449
rect 243358 7375 243414 7384
rect 243372 7154 243400 7375
rect 243634 7168 243690 7177
rect 243372 7126 243634 7154
rect 243634 7103 243690 7112
rect 243542 3768 243598 3777
rect 243542 3703 243598 3712
rect 243556 3097 243584 3703
rect 243542 3088 243598 3097
rect 243542 3023 243598 3032
rect 246408 480 246436 79591
rect 260654 10568 260710 10577
rect 260654 10503 260710 10512
rect 249982 8120 250038 8129
rect 249982 8055 250038 8064
rect 248326 3768 248382 3777
rect 248326 3703 248382 3712
rect 248340 2961 248368 3703
rect 248326 2952 248382 2961
rect 248326 2887 248382 2896
rect 249996 480 250024 8055
rect 256700 7880 256752 7886
rect 256700 7822 256752 7828
rect 253204 7744 253256 7750
rect 253204 7686 253256 7692
rect 251088 7608 251140 7614
rect 251088 7550 251140 7556
rect 251100 7449 251128 7550
rect 251086 7440 251142 7449
rect 251086 7375 251142 7384
rect 253216 7041 253244 7686
rect 256712 7449 256740 7822
rect 256698 7440 256754 7449
rect 256698 7375 256754 7384
rect 257066 7440 257122 7449
rect 257066 7375 257122 7384
rect 253478 7304 253534 7313
rect 253478 7239 253534 7248
rect 253202 7032 253258 7041
rect 253202 6967 253258 6976
rect 253492 480 253520 7239
rect 257080 480 257108 7375
rect 260668 480 260696 10503
rect 263782 7304 263838 7313
rect 263782 7239 263838 7248
rect 263796 7154 263824 7239
rect 264058 7168 264114 7177
rect 263796 7126 264058 7154
rect 264058 7103 264114 7112
rect 264164 480 264192 120119
rect 265622 7304 265678 7313
rect 265622 7239 265678 7248
rect 265636 7041 265664 7239
rect 265622 7032 265678 7041
rect 265622 6967 265678 6976
rect 267752 480 267780 120527
rect 271234 120456 271290 120465
rect 271234 120391 271290 120400
rect 271248 480 271276 120391
rect 274822 120320 274878 120329
rect 274822 120255 274878 120264
rect 273166 7168 273222 7177
rect 273442 7168 273498 7177
rect 273222 7126 273442 7154
rect 273166 7103 273222 7112
rect 273442 7103 273498 7112
rect 274836 480 274864 120255
rect 304552 118660 304580 120527
rect 313646 120456 313702 120465
rect 313646 120391 313702 120400
rect 313660 118660 313688 120391
rect 322754 120320 322810 120329
rect 322754 120255 322810 120264
rect 322768 118660 322796 120255
rect 331862 120184 331918 120193
rect 331862 120119 331918 120128
rect 331876 118660 331904 120119
rect 339774 115560 339830 115569
rect 339774 115495 339830 115504
rect 338118 114608 338174 114617
rect 338118 114543 338174 114552
rect 337474 112704 337530 112713
rect 337474 112639 337530 112648
rect 336002 108352 336058 108361
rect 336002 108287 336058 108296
rect 302436 78062 302464 80036
rect 306944 78441 306972 80036
rect 306930 78432 306986 78441
rect 306930 78367 306986 78376
rect 305644 78124 305696 78130
rect 305644 78066 305696 78072
rect 302424 78056 302476 78062
rect 302424 77998 302476 78004
rect 300122 77752 300178 77761
rect 300122 77687 300178 77696
rect 300136 9081 300164 77687
rect 300122 9072 300178 9081
rect 300122 9007 300178 9016
rect 303158 9072 303214 9081
rect 303158 9007 303214 9016
rect 299662 8936 299718 8945
rect 299662 8871 299718 8880
rect 292578 8800 292634 8809
rect 292578 8735 292634 8744
rect 278318 8664 278374 8673
rect 278318 8599 278374 8608
rect 275282 7304 275338 7313
rect 275282 7239 275338 7248
rect 275296 7041 275324 7239
rect 275282 7032 275338 7041
rect 275282 6967 275338 6976
rect 278332 480 278360 8599
rect 284942 7304 284998 7313
rect 284942 7239 284998 7248
rect 282918 7168 282974 7177
rect 283194 7168 283250 7177
rect 282974 7126 283194 7154
rect 282918 7103 282974 7112
rect 283194 7103 283250 7112
rect 284956 7041 284984 7239
rect 284942 7032 284998 7041
rect 284942 6967 284998 6976
rect 285588 5500 285640 5506
rect 285588 5442 285640 5448
rect 285402 5128 285458 5137
rect 285402 5063 285458 5072
rect 281906 4992 281962 5001
rect 281906 4927 281962 4936
rect 281920 480 281948 4927
rect 285416 480 285444 5063
rect 285600 4321 285628 5442
rect 288440 5432 288492 5438
rect 288440 5374 288492 5380
rect 288990 5400 289046 5409
rect 288452 4457 288480 5374
rect 288990 5335 289046 5344
rect 288438 4448 288494 4457
rect 288438 4383 288494 4392
rect 285586 4312 285642 4321
rect 285586 4247 285642 4256
rect 289004 480 289032 5335
rect 292592 480 292620 8735
rect 294602 7304 294658 7313
rect 294602 7239 294658 7248
rect 292670 7168 292726 7177
rect 292946 7168 293002 7177
rect 292726 7126 292946 7154
rect 292670 7103 292726 7112
rect 292946 7103 293002 7112
rect 294616 7041 294644 7239
rect 294602 7032 294658 7041
rect 294602 6967 294658 6976
rect 296074 2952 296130 2961
rect 296074 2887 296130 2896
rect 296088 480 296116 2887
rect 299676 480 299704 8871
rect 303172 480 303200 9007
rect 305656 5506 305684 78066
rect 307024 78056 307076 78062
rect 307024 77998 307076 78004
rect 305644 5500 305696 5506
rect 305644 5442 305696 5448
rect 307036 5438 307064 77998
rect 310242 9208 310298 9217
rect 310242 9143 310298 9152
rect 307668 5500 307720 5506
rect 307668 5442 307720 5448
rect 307024 5432 307076 5438
rect 307024 5374 307076 5380
rect 306746 4720 306802 4729
rect 306746 4655 306802 4664
rect 306760 480 306788 4655
rect 307680 4185 307708 5442
rect 307666 4176 307722 4185
rect 307666 4111 307722 4120
rect 310256 480 310284 9143
rect 311452 4865 311480 80036
rect 315960 78305 315988 80036
rect 315946 78296 316002 78305
rect 315946 78231 316002 78240
rect 320468 78169 320496 80036
rect 324976 78577 325004 80036
rect 329484 78674 329512 80036
rect 329472 78668 329524 78674
rect 329472 78610 329524 78616
rect 324962 78568 325018 78577
rect 324962 78503 325018 78512
rect 320824 78192 320876 78198
rect 320454 78160 320510 78169
rect 320824 78134 320876 78140
rect 327998 78160 328054 78169
rect 320454 78095 320510 78104
rect 320836 9654 320864 78134
rect 327998 78095 328054 78104
rect 313280 9648 313332 9654
rect 313280 9590 313332 9596
rect 320824 9648 320876 9654
rect 325608 9648 325660 9654
rect 320824 9590 320876 9596
rect 320914 9616 320970 9625
rect 313292 8537 313320 9590
rect 320732 9580 320784 9586
rect 325608 9590 325660 9596
rect 320914 9551 320970 9560
rect 320732 9522 320784 9528
rect 317328 9512 317380 9518
rect 317234 9480 317290 9489
rect 317328 9454 317380 9460
rect 317234 9415 317290 9424
rect 313830 9344 313886 9353
rect 313830 9279 313886 9288
rect 313278 8528 313334 8537
rect 313278 8463 313334 8472
rect 311438 4856 311494 4865
rect 311438 4791 311494 4800
rect 313844 480 313872 9279
rect 317248 6914 317276 9415
rect 317340 8401 317368 9454
rect 320744 8673 320772 9522
rect 320730 8664 320786 8673
rect 320730 8599 320786 8608
rect 317326 8392 317382 8401
rect 317326 8327 317382 8336
rect 317248 6886 317368 6914
rect 317340 480 317368 6886
rect 320928 480 320956 9551
rect 325620 8809 325648 9590
rect 325606 8800 325662 8809
rect 325606 8735 325662 8744
rect 324410 8664 324466 8673
rect 324410 8599 324466 8608
rect 323582 7304 323638 7313
rect 323582 7239 323638 7248
rect 321558 7168 321614 7177
rect 321834 7168 321890 7177
rect 321614 7126 321834 7154
rect 321558 7103 321614 7112
rect 321834 7103 321890 7112
rect 323596 7041 323624 7239
rect 323582 7032 323638 7041
rect 323582 6967 323638 6976
rect 324424 480 324452 8599
rect 328012 480 328040 78095
rect 333992 77994 334020 80036
rect 335082 78296 335138 78305
rect 335082 78231 335138 78240
rect 333980 77988 334032 77994
rect 333980 77930 334032 77936
rect 331586 4856 331642 4865
rect 331586 4791 331642 4800
rect 331600 480 331628 4791
rect 335096 480 335124 78231
rect 335542 8256 335598 8265
rect 335542 8191 335598 8200
rect 335556 7886 335584 8191
rect 335726 8120 335782 8129
rect 335726 8055 335782 8064
rect 335544 7880 335596 7886
rect 335544 7822 335596 7828
rect 335740 7750 335768 8055
rect 335728 7744 335780 7750
rect 335728 7686 335780 7692
rect 336016 6914 336044 108287
rect 336830 106992 336886 107001
rect 336830 106927 336886 106936
rect 336738 105088 336794 105097
rect 336738 105023 336794 105032
rect 336094 96928 336150 96937
rect 336094 96863 336150 96872
rect 336108 8378 336136 96863
rect 336278 89584 336334 89593
rect 336278 89519 336334 89528
rect 336186 88360 336242 88369
rect 336186 88295 336242 88304
rect 336200 9518 336228 88295
rect 336188 9512 336240 9518
rect 336188 9454 336240 9460
rect 336108 8350 336228 8378
rect 336094 8256 336150 8265
rect 336094 8191 336150 8200
rect 336108 7614 336136 8191
rect 336096 7608 336148 7614
rect 336096 7550 336148 7556
rect 336200 7449 336228 8350
rect 336292 7585 336320 89519
rect 336370 87272 336426 87281
rect 336370 87207 336426 87216
rect 336278 7576 336334 7585
rect 336278 7511 336334 7520
rect 336186 7440 336242 7449
rect 336186 7375 336242 7384
rect 336384 7177 336412 87207
rect 336554 81560 336610 81569
rect 336554 81495 336610 81504
rect 336568 80102 336596 81495
rect 336752 80186 336780 105023
rect 336660 80158 336780 80186
rect 336556 80096 336608 80102
rect 336660 80073 336688 80158
rect 336740 80096 336792 80102
rect 336556 80038 336608 80044
rect 336646 80064 336702 80073
rect 336740 80038 336792 80044
rect 336646 79999 336702 80008
rect 336752 77625 336780 80038
rect 336738 77616 336794 77625
rect 336738 77551 336794 77560
rect 336844 10577 336872 106927
rect 336922 103184 336978 103193
rect 336922 103119 336978 103128
rect 336830 10568 336886 10577
rect 336830 10503 336886 10512
rect 336370 7168 336426 7177
rect 336370 7103 336426 7112
rect 335924 6886 336044 6914
rect 335924 5506 335952 6886
rect 336936 6089 336964 103119
rect 337382 101280 337438 101289
rect 337382 101215 337438 101224
rect 337014 95568 337070 95577
rect 337014 95503 337070 95512
rect 337028 7993 337056 95503
rect 337106 93664 337162 93673
rect 337106 93599 337162 93608
rect 337014 7984 337070 7993
rect 337014 7919 337070 7928
rect 337120 6905 337148 93599
rect 337198 91760 337254 91769
rect 337198 91695 337254 91704
rect 337106 6896 337162 6905
rect 337106 6831 337162 6840
rect 337212 6633 337240 91695
rect 337290 86048 337346 86057
rect 337290 85983 337346 85992
rect 337304 7857 337332 85983
rect 337396 80306 337424 101215
rect 337488 89714 337516 112639
rect 337488 89686 337700 89714
rect 337384 80300 337436 80306
rect 337384 80242 337436 80248
rect 337384 80096 337436 80102
rect 337672 80054 337700 89686
rect 337384 80038 337436 80044
rect 337396 22681 337424 80038
rect 337488 80026 337700 80054
rect 337382 22672 337438 22681
rect 337382 22607 337438 22616
rect 337290 7848 337346 7857
rect 337290 7783 337346 7792
rect 337488 7721 337516 80026
rect 338132 8265 338160 114543
rect 339498 113656 339554 113665
rect 339498 113591 339554 113600
rect 338302 104136 338358 104145
rect 338302 104071 338358 104080
rect 338210 102232 338266 102241
rect 338210 102167 338266 102176
rect 338118 8256 338174 8265
rect 338118 8191 338174 8200
rect 337474 7712 337530 7721
rect 337474 7647 337530 7656
rect 337198 6624 337254 6633
rect 337198 6559 337254 6568
rect 338224 6225 338252 102167
rect 338316 85270 338344 104071
rect 338854 96520 338910 96529
rect 338854 96455 338910 96464
rect 338486 94616 338542 94625
rect 338486 94551 338542 94560
rect 338394 92712 338450 92721
rect 338394 92647 338450 92656
rect 338304 85264 338356 85270
rect 338304 85206 338356 85212
rect 338302 83192 338358 83201
rect 338302 83127 338358 83136
rect 338316 79393 338344 83127
rect 338302 79384 338358 79393
rect 338302 79319 338358 79328
rect 338408 6914 338436 92647
rect 338316 6886 338436 6914
rect 338210 6216 338266 6225
rect 338210 6151 338266 6160
rect 336922 6080 336978 6089
rect 336922 6015 336978 6024
rect 335912 5500 335964 5506
rect 335912 5442 335964 5448
rect 336648 4820 336700 4826
rect 336648 4762 336700 4768
rect 335174 4176 335230 4185
rect 335174 4111 335230 4120
rect 335188 3777 335216 4111
rect 335174 3768 335230 3777
rect 335174 3703 335230 3712
rect 336660 3534 336688 4762
rect 338316 3777 338344 6886
rect 338500 6497 338528 94551
rect 338578 90808 338634 90817
rect 338578 90743 338634 90752
rect 338592 6866 338620 90743
rect 338762 87000 338818 87009
rect 338762 86935 338818 86944
rect 338672 85264 338724 85270
rect 338672 85206 338724 85212
rect 338684 81161 338712 85206
rect 338670 81152 338726 81161
rect 338670 81087 338726 81096
rect 338776 80054 338804 86935
rect 338684 80026 338804 80054
rect 338580 6860 338632 6866
rect 338580 6802 338632 6808
rect 338486 6488 338542 6497
rect 338486 6423 338542 6432
rect 338684 5273 338712 80026
rect 338868 79490 338896 96455
rect 338946 85096 339002 85105
rect 338946 85031 339002 85040
rect 338856 79484 338908 79490
rect 338856 79426 338908 79432
rect 338960 79370 338988 85031
rect 338776 79342 338988 79370
rect 338776 6361 338804 79342
rect 338856 79280 338908 79286
rect 338856 79222 338908 79228
rect 338762 6352 338818 6361
rect 338762 6287 338818 6296
rect 338868 5545 338896 79222
rect 338854 5536 338910 5545
rect 338854 5471 338910 5480
rect 338670 5264 338726 5273
rect 338670 5199 338726 5208
rect 338486 4040 338542 4049
rect 338486 3975 338542 3984
rect 338670 4040 338726 4049
rect 338670 3975 338726 3984
rect 338500 3777 338528 3975
rect 338302 3768 338358 3777
rect 338302 3703 338358 3712
rect 338486 3768 338542 3777
rect 338486 3703 338542 3712
rect 336648 3528 336700 3534
rect 336648 3470 336700 3476
rect 338684 480 338712 3975
rect 339512 3777 339540 113591
rect 339590 100328 339646 100337
rect 339590 100263 339646 100272
rect 339498 3768 339554 3777
rect 339498 3703 339554 3712
rect 339604 3466 339632 100263
rect 339682 84144 339738 84153
rect 339682 84079 339738 84088
rect 339592 3460 339644 3466
rect 339592 3402 339644 3408
rect 339696 3233 339724 84079
rect 339788 79529 339816 115495
rect 398102 107808 398158 107817
rect 398102 107743 398158 107752
rect 398116 79966 398144 107743
rect 398104 79960 398156 79966
rect 398104 79902 398156 79908
rect 339774 79520 339830 79529
rect 339774 79455 339830 79464
rect 400968 78198 400996 80036
rect 400956 78192 401008 78198
rect 400956 78134 401008 78140
rect 402532 4826 402560 80036
rect 403622 78432 403678 78441
rect 403622 78367 403678 78376
rect 402520 4820 402572 4826
rect 402520 4762 402572 4768
rect 344926 4176 344982 4185
rect 344926 4111 344982 4120
rect 344940 3777 344968 4111
rect 349710 4040 349766 4049
rect 349710 3975 349766 3984
rect 356150 4040 356206 4049
rect 356150 3975 356206 3984
rect 356334 4040 356390 4049
rect 356334 3975 356390 3984
rect 398102 4040 398158 4049
rect 398102 3975 398158 3984
rect 398286 4040 398342 4049
rect 398286 3975 398342 3984
rect 349724 3890 349752 3975
rect 349986 3904 350042 3913
rect 349724 3862 349986 3890
rect 349986 3839 350042 3848
rect 344926 3768 344982 3777
rect 344926 3703 344982 3712
rect 356164 3233 356192 3975
rect 339682 3224 339738 3233
rect 339682 3159 339738 3168
rect 356150 3224 356206 3233
rect 356150 3159 356206 3168
rect 356348 480 356376 3975
rect 398116 3233 398144 3975
rect 398102 3224 398158 3233
rect 398102 3159 398158 3168
rect 398300 3097 398328 3975
rect 403636 3233 403664 78367
rect 404096 4078 404124 80036
rect 405660 4146 405688 80036
rect 405648 4140 405700 4146
rect 405648 4082 405700 4088
rect 404084 4072 404136 4078
rect 404084 4014 404136 4020
rect 407224 4010 407252 80036
rect 408788 78130 408816 80036
rect 408776 78124 408828 78130
rect 408776 78066 408828 78072
rect 407762 77888 407818 77897
rect 407762 77823 407818 77832
rect 407776 77489 407804 77823
rect 407762 77480 407818 77489
rect 407762 77415 407818 77424
rect 410352 77353 410380 80036
rect 411916 78062 411944 80036
rect 411904 78056 411956 78062
rect 411904 77998 411956 78004
rect 413480 77897 413508 80036
rect 414662 78568 414718 78577
rect 414662 78503 414718 78512
rect 413466 77888 413522 77897
rect 413466 77823 413522 77832
rect 411994 77616 412050 77625
rect 411994 77551 412050 77560
rect 410338 77344 410394 77353
rect 410338 77279 410394 77288
rect 407212 4004 407264 4010
rect 407212 3946 407264 3952
rect 412008 3641 412036 77551
rect 414676 4049 414704 78503
rect 415044 77489 415072 80036
rect 416608 77625 416636 80036
rect 418172 78033 418200 80036
rect 418158 78024 418214 78033
rect 418158 77959 418214 77968
rect 416594 77616 416650 77625
rect 416594 77551 416650 77560
rect 415030 77480 415086 77489
rect 415030 77415 415086 77424
rect 414662 4040 414718 4049
rect 414662 3975 414718 3984
rect 411994 3632 412050 3641
rect 411994 3567 412050 3576
rect 419736 3505 419764 80036
rect 421300 77761 421328 80036
rect 422864 78577 422892 80036
rect 422850 78568 422906 78577
rect 422850 78503 422906 78512
rect 421286 77752 421342 77761
rect 421286 77687 421342 77696
rect 424428 9586 424456 80036
rect 424416 9580 424468 9586
rect 424416 9522 424468 9528
rect 425992 5001 426020 80036
rect 427556 5137 427584 80036
rect 429120 5409 429148 80036
rect 430684 9654 430712 80036
rect 432248 78577 432276 80036
rect 432234 78568 432290 78577
rect 432234 78503 432290 78512
rect 430672 9648 430724 9654
rect 430672 9590 430724 9596
rect 433812 8945 433840 80036
rect 435376 9081 435404 80036
rect 435362 9072 435418 9081
rect 435362 9007 435418 9016
rect 433798 8936 433854 8945
rect 433798 8871 433854 8880
rect 429106 5400 429162 5409
rect 429106 5335 429162 5344
rect 427542 5128 427598 5137
rect 427542 5063 427598 5072
rect 425978 4992 426034 5001
rect 425978 4927 426034 4936
rect 436940 4729 436968 80036
rect 438504 9217 438532 80036
rect 440068 9353 440096 80036
rect 441632 9489 441660 80036
rect 443196 9625 443224 80036
rect 443182 9616 443238 9625
rect 443182 9551 443238 9560
rect 441618 9480 441674 9489
rect 441618 9415 441674 9424
rect 440054 9344 440110 9353
rect 440054 9279 440110 9288
rect 438490 9208 438546 9217
rect 438490 9143 438546 9152
rect 444760 8673 444788 80036
rect 446324 78169 446352 80036
rect 446310 78160 446366 78169
rect 446310 78095 446366 78104
rect 444746 8664 444802 8673
rect 444746 8599 444802 8608
rect 447888 4865 447916 80036
rect 449452 78305 449480 80036
rect 449438 78296 449494 78305
rect 449438 78231 449494 78240
rect 447874 4856 447930 4865
rect 447874 4791 447930 4800
rect 436926 4720 436982 4729
rect 436926 4655 436982 4664
rect 451016 3913 451044 80036
rect 452580 78441 452608 80036
rect 452566 78432 452622 78441
rect 452566 78367 452622 78376
rect 451002 3904 451058 3913
rect 451002 3839 451058 3848
rect 419722 3496 419778 3505
rect 419722 3431 419778 3440
rect 403622 3224 403678 3233
rect 403622 3159 403678 3168
rect 398286 3088 398342 3097
rect 398286 3023 398342 3032
rect 97418 326 97856 354
rect 97418 -960 97530 326
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 348790 700440 348846 700496
rect 109038 700304 109094 700360
rect 104714 697176 104770 697232
rect 100390 644000 100446 644056
rect 96066 590960 96122 591016
rect 91742 537784 91798 537840
rect 87418 484608 87474 484664
rect 83094 298696 83150 298752
rect 152278 630808 152334 630864
rect 147954 577632 148010 577688
rect 143630 524456 143686 524512
rect 139306 471416 139362 471472
rect 118054 192616 118110 192672
rect 113638 192480 113694 192536
rect 397458 192616 397514 192672
rect 527178 700304 527234 700360
rect 462318 192480 462374 192536
rect 191838 186496 191894 186552
rect 190458 164600 190514 164656
rect 189998 135768 190054 135824
rect 189354 123392 189410 123448
rect 4066 77968 4122 78024
rect 1674 6568 1730 6624
rect 570 5616 626 5672
rect 2870 3032 2926 3088
rect 5262 77832 5318 77888
rect 41878 77424 41934 77480
rect 18234 77288 18290 77344
rect 7654 6704 7710 6760
rect 6458 3712 6514 3768
rect 13542 6160 13598 6216
rect 9954 5752 10010 5808
rect 8758 4120 8814 4176
rect 12346 2760 12402 2816
rect 17038 4800 17094 4856
rect 14738 2896 14794 2952
rect 32402 11056 32458 11112
rect 31298 10240 31354 10296
rect 23018 9696 23074 9752
rect 21822 4936 21878 4992
rect 19430 2760 19486 2816
rect 30102 5208 30158 5264
rect 26514 5072 26570 5128
rect 24214 3576 24270 3632
rect 27710 3440 27766 3496
rect 28906 3304 28962 3360
rect 38382 10512 38438 10568
rect 34794 10376 34850 10432
rect 33598 5344 33654 5400
rect 37186 5480 37242 5536
rect 35990 3848 36046 3904
rect 40774 4664 40830 4720
rect 40682 4120 40738 4176
rect 40682 3984 40738 4040
rect 40682 3576 40738 3632
rect 39578 3440 39634 3496
rect 67914 12960 67970 13016
rect 64326 12008 64382 12064
rect 60830 11872 60886 11928
rect 53746 11736 53802 11792
rect 50158 11600 50214 11656
rect 46662 11192 46718 11248
rect 45466 10648 45522 10704
rect 44270 9152 44326 9208
rect 43074 3168 43130 3224
rect 47858 6840 47914 6896
rect 51354 7384 51410 7440
rect 52550 6296 52606 6352
rect 56046 8472 56102 8528
rect 54942 7928 54998 7984
rect 59634 8336 59690 8392
rect 58438 7112 58494 7168
rect 57242 3168 57298 3224
rect 63222 8608 63278 8664
rect 62026 6976 62082 7032
rect 65522 7248 65578 7304
rect 66718 3168 66774 3224
rect 74998 12280 75054 12336
rect 71502 12144 71558 12200
rect 70306 8880 70362 8936
rect 69110 3168 69166 3224
rect 72606 7520 72662 7576
rect 73802 6432 73858 6488
rect 73158 5616 73214 5672
rect 78494 11464 78550 11520
rect 75826 11056 75882 11112
rect 77390 9016 77446 9072
rect 77206 5752 77262 5808
rect 76194 5616 76250 5672
rect 78586 11192 78642 11248
rect 80886 10784 80942 10840
rect 79690 7656 79746 7712
rect 83094 7792 83150 7848
rect 83278 7792 83334 7848
rect 82818 7384 82874 7440
rect 83094 7384 83150 7440
rect 82082 3168 82138 3224
rect 81438 3032 81494 3088
rect 84842 77968 84898 78024
rect 86406 77832 86462 77888
rect 84474 10920 84530 10976
rect 83370 6568 83426 6624
rect 87970 10104 88026 10160
rect 86866 7928 86922 7984
rect 87050 7928 87106 7984
rect 88246 9696 88302 9752
rect 91558 78240 91614 78296
rect 91098 77288 91154 77344
rect 90362 9288 90418 9344
rect 89626 6704 89682 6760
rect 89166 6568 89222 6624
rect 88062 3576 88118 3632
rect 88982 3576 89038 3632
rect 88982 3168 89038 3224
rect 89718 3848 89774 3904
rect 93950 9424 94006 9480
rect 92754 6704 92810 6760
rect 92662 4800 92718 4856
rect 95146 8472 95202 8528
rect 98642 77832 98698 77888
rect 97814 9560 97870 9616
rect 97446 5208 97502 5264
rect 95882 5072 95938 5128
rect 94318 4936 94374 4992
rect 95146 3712 95202 3768
rect 96250 3712 96306 3768
rect 97906 8608 97962 8664
rect 98550 7384 98606 7440
rect 98826 7112 98882 7168
rect 101034 8744 101090 8800
rect 100758 8336 100814 8392
rect 100574 5480 100630 5536
rect 99010 5344 99066 5400
rect 99838 3984 99894 4040
rect 102230 77968 102286 78024
rect 102138 4664 102194 4720
rect 102138 2896 102194 2952
rect 103702 9152 103758 9208
rect 104530 8064 104586 8120
rect 103334 3168 103390 3224
rect 104806 7384 104862 7440
rect 105726 78512 105782 78568
rect 105266 6840 105322 6896
rect 108118 8200 108174 8256
rect 107658 6976 107714 7032
rect 106922 6840 106978 6896
rect 112810 77696 112866 77752
rect 110418 7248 110474 7304
rect 111614 7384 111670 7440
rect 116122 78104 116178 78160
rect 116122 77560 116178 77616
rect 114650 77288 114706 77344
rect 116398 77560 116454 77616
rect 116214 7520 116270 7576
rect 115202 4800 115258 4856
rect 114006 2896 114062 2952
rect 117226 77424 117282 77480
rect 118698 78104 118754 78160
rect 119894 77424 119950 77480
rect 119342 7656 119398 7712
rect 117778 6024 117834 6080
rect 118790 5344 118846 5400
rect 117594 4936 117650 4992
rect 123482 77288 123538 77344
rect 122470 7928 122526 7984
rect 120906 7792 120962 7848
rect 122286 5480 122342 5536
rect 121090 5072 121146 5128
rect 124126 78240 124182 78296
rect 127162 9560 127218 9616
rect 125598 9424 125654 9480
rect 124034 9288 124090 9344
rect 128726 8744 128782 8800
rect 131854 8200 131910 8256
rect 130290 8064 130346 8120
rect 133418 7384 133474 7440
rect 124678 5208 124734 5264
rect 138110 5480 138166 5536
rect 144918 77852 144974 77888
rect 144918 77832 144920 77852
rect 144920 77832 144972 77852
rect 144972 77832 144974 77852
rect 145838 77832 145894 77888
rect 146022 77852 146078 77888
rect 146022 77832 146024 77852
rect 146024 77832 146076 77852
rect 146076 77832 146078 77852
rect 153750 10648 153806 10704
rect 150622 10512 150678 10568
rect 149058 10376 149114 10432
rect 147494 10240 147550 10296
rect 154210 7656 154266 7712
rect 141238 6160 141294 6216
rect 136546 5344 136602 5400
rect 134982 4800 135038 4856
rect 155406 8336 155462 8392
rect 158902 10240 158958 10296
rect 156878 6296 156934 6352
rect 157798 5616 157854 5672
rect 156602 5344 156658 5400
rect 163042 78104 163098 78160
rect 164882 10376 164938 10432
rect 164698 8880 164754 8936
rect 162490 6976 162546 7032
rect 160098 6296 160154 6352
rect 163686 4800 163742 4856
rect 166078 7112 166134 7168
rect 168378 79328 168434 79384
rect 167826 9016 167882 9072
rect 166262 6432 166318 6488
rect 167182 5480 167238 5536
rect 170954 10920 171010 10976
rect 169390 10784 169446 10840
rect 172518 10104 172574 10160
rect 169574 7520 169630 7576
rect 177118 77968 177174 78024
rect 175554 77832 175610 77888
rect 180246 78512 180302 78568
rect 178682 78376 178738 78432
rect 179234 78376 179290 78432
rect 178958 78104 179014 78160
rect 175462 6160 175518 6216
rect 174542 5344 174598 5400
rect 170770 4664 170826 4720
rect 172978 4256 173034 4312
rect 171966 3032 172022 3088
rect 174266 4120 174322 4176
rect 172978 3848 173034 3904
rect 173162 3848 173218 3904
rect 173622 3848 173678 3904
rect 172426 2760 172482 2816
rect 173622 3032 173678 3088
rect 176658 4392 176714 4448
rect 180062 78240 180118 78296
rect 179234 6296 179290 6352
rect 179050 5752 179106 5808
rect 178958 4664 179014 4720
rect 180246 7384 180302 7440
rect 180062 5480 180118 5536
rect 181074 7384 181130 7440
rect 180798 7248 180854 7304
rect 183374 77696 183430 77752
rect 184938 77560 184994 77616
rect 186502 77424 186558 77480
rect 188066 77288 188122 77344
rect 189446 120264 189502 120320
rect 189354 11736 189410 11792
rect 189538 110880 189594 110936
rect 189446 11600 189502 11656
rect 183742 8472 183798 8528
rect 182546 6296 182602 6352
rect 185582 6432 185638 6488
rect 185582 6024 185638 6080
rect 186134 6432 186190 6488
rect 185674 5616 185730 5672
rect 185582 3440 185638 3496
rect 185030 3304 185086 3360
rect 185582 3032 185638 3088
rect 185030 2896 185086 2952
rect 189630 101496 189686 101552
rect 189538 3440 189594 3496
rect 189906 95240 189962 95296
rect 189814 88848 189870 88904
rect 189722 80552 189778 80608
rect 189722 7656 189778 7712
rect 189998 12960 190054 13016
rect 190550 161472 190606 161528
rect 190458 3984 190514 4040
rect 190642 152088 190698 152144
rect 190734 145832 190790 145888
rect 190826 142704 190882 142760
rect 190918 139576 190974 139632
rect 190826 12280 190882 12336
rect 191010 133320 191066 133376
rect 190918 12144 190974 12200
rect 191102 130192 191158 130248
rect 191010 12008 191066 12064
rect 191194 117680 191250 117736
rect 191286 105168 191342 105224
rect 191102 11872 191158 11928
rect 190734 11464 190790 11520
rect 191930 183368 191986 183424
rect 191838 5208 191894 5264
rect 192022 180240 192078 180296
rect 191930 5072 191986 5128
rect 192114 173984 192170 174040
rect 192206 170856 192262 170912
rect 192298 167728 192354 167784
rect 192206 6840 192262 6896
rect 192114 5480 192170 5536
rect 192022 4936 192078 4992
rect 190826 3984 190882 4040
rect 190550 3712 190606 3768
rect 189722 3440 189778 3496
rect 189630 2896 189686 2952
rect 192390 158344 192446 158400
rect 192482 155216 192538 155272
rect 192390 6568 192446 6624
rect 192574 148960 192630 149016
rect 192482 6024 192538 6080
rect 192298 3168 192354 3224
rect 267738 120536 267794 120592
rect 304538 120536 304594 120592
rect 264150 120128 264206 120184
rect 192666 108296 192722 108352
rect 193862 80688 193918 80744
rect 193218 3984 193274 4040
rect 192574 3032 192630 3088
rect 190826 2896 190882 2952
rect 246394 79600 246450 79656
rect 207386 79464 207442 79520
rect 200302 5480 200358 5536
rect 196806 5208 196862 5264
rect 193862 3440 193918 3496
rect 194414 3032 194470 3088
rect 197910 2760 197966 2816
rect 201498 4256 201554 4312
rect 205086 3712 205142 3768
rect 203890 3168 203946 3224
rect 222750 77968 222806 78024
rect 215666 77832 215722 77888
rect 210974 77560 211030 77616
rect 208582 4392 208638 4448
rect 214470 6568 214526 6624
rect 212170 3304 212226 3360
rect 218058 22616 218114 22672
rect 222106 6976 222162 7032
rect 221554 6704 221610 6760
rect 219254 3576 219310 3632
rect 229834 9016 229890 9072
rect 222842 7404 222898 7440
rect 222842 7384 222844 7404
rect 222844 7384 222896 7404
rect 222896 7384 222898 7404
rect 228730 6840 228786 6896
rect 226338 3440 226394 3496
rect 225142 3168 225198 3224
rect 224958 2896 225014 2952
rect 226430 3032 226486 3088
rect 242898 7928 242954 7984
rect 239310 7792 239366 7848
rect 235814 7656 235870 7712
rect 232226 6024 232282 6080
rect 233238 3712 233294 3768
rect 233422 3712 233478 3768
rect 233238 2896 233294 2952
rect 233882 2760 233938 2816
rect 243358 7384 243414 7440
rect 243634 7112 243690 7168
rect 243542 3712 243598 3768
rect 243542 3032 243598 3088
rect 260654 10512 260710 10568
rect 249982 8064 250038 8120
rect 248326 3712 248382 3768
rect 248326 2896 248382 2952
rect 251086 7384 251142 7440
rect 256698 7384 256754 7440
rect 257066 7384 257122 7440
rect 253478 7248 253534 7304
rect 253202 6976 253258 7032
rect 263782 7248 263838 7304
rect 264058 7112 264114 7168
rect 265622 7248 265678 7304
rect 265622 6976 265678 7032
rect 271234 120400 271290 120456
rect 274822 120264 274878 120320
rect 273166 7112 273222 7168
rect 273442 7112 273498 7168
rect 313646 120400 313702 120456
rect 322754 120264 322810 120320
rect 331862 120128 331918 120184
rect 339774 115504 339830 115560
rect 338118 114552 338174 114608
rect 337474 112648 337530 112704
rect 336002 108296 336058 108352
rect 306930 78376 306986 78432
rect 300122 77696 300178 77752
rect 300122 9016 300178 9072
rect 303158 9016 303214 9072
rect 299662 8880 299718 8936
rect 292578 8744 292634 8800
rect 278318 8608 278374 8664
rect 275282 7248 275338 7304
rect 275282 6976 275338 7032
rect 284942 7248 284998 7304
rect 282918 7112 282974 7168
rect 283194 7112 283250 7168
rect 284942 6976 284998 7032
rect 285402 5072 285458 5128
rect 281906 4936 281962 4992
rect 288990 5344 289046 5400
rect 288438 4392 288494 4448
rect 285586 4256 285642 4312
rect 294602 7248 294658 7304
rect 292670 7112 292726 7168
rect 292946 7112 293002 7168
rect 294602 6976 294658 7032
rect 296074 2896 296130 2952
rect 310242 9152 310298 9208
rect 306746 4664 306802 4720
rect 307666 4120 307722 4176
rect 315946 78240 316002 78296
rect 324962 78512 325018 78568
rect 320454 78104 320510 78160
rect 327998 78104 328054 78160
rect 320914 9560 320970 9616
rect 317234 9424 317290 9480
rect 313830 9288 313886 9344
rect 313278 8472 313334 8528
rect 311438 4800 311494 4856
rect 320730 8608 320786 8664
rect 317326 8336 317382 8392
rect 325606 8744 325662 8800
rect 324410 8608 324466 8664
rect 323582 7248 323638 7304
rect 321558 7112 321614 7168
rect 321834 7112 321890 7168
rect 323582 6976 323638 7032
rect 335082 78240 335138 78296
rect 331586 4800 331642 4856
rect 335542 8200 335598 8256
rect 335726 8064 335782 8120
rect 336830 106936 336886 106992
rect 336738 105032 336794 105088
rect 336094 96872 336150 96928
rect 336278 89528 336334 89584
rect 336186 88304 336242 88360
rect 336094 8200 336150 8256
rect 336370 87216 336426 87272
rect 336278 7520 336334 7576
rect 336186 7384 336242 7440
rect 336554 81504 336610 81560
rect 336646 80008 336702 80064
rect 336738 77560 336794 77616
rect 336922 103128 336978 103184
rect 336830 10512 336886 10568
rect 336370 7112 336426 7168
rect 337382 101224 337438 101280
rect 337014 95512 337070 95568
rect 337106 93608 337162 93664
rect 337014 7928 337070 7984
rect 337198 91704 337254 91760
rect 337106 6840 337162 6896
rect 337290 85992 337346 86048
rect 337382 22616 337438 22672
rect 337290 7792 337346 7848
rect 339498 113600 339554 113656
rect 338302 104080 338358 104136
rect 338210 102176 338266 102232
rect 338118 8200 338174 8256
rect 337474 7656 337530 7712
rect 337198 6568 337254 6624
rect 338854 96464 338910 96520
rect 338486 94560 338542 94616
rect 338394 92656 338450 92712
rect 338302 83136 338358 83192
rect 338302 79328 338358 79384
rect 338210 6160 338266 6216
rect 336922 6024 336978 6080
rect 335174 4120 335230 4176
rect 335174 3712 335230 3768
rect 338578 90752 338634 90808
rect 338762 86944 338818 87000
rect 338670 81096 338726 81152
rect 338486 6432 338542 6488
rect 338946 85040 339002 85096
rect 338762 6296 338818 6352
rect 338854 5480 338910 5536
rect 338670 5208 338726 5264
rect 338486 3984 338542 4040
rect 338670 3984 338726 4040
rect 338302 3712 338358 3768
rect 338486 3712 338542 3768
rect 339590 100272 339646 100328
rect 339498 3712 339554 3768
rect 339682 84088 339738 84144
rect 398102 107752 398158 107808
rect 339774 79464 339830 79520
rect 403622 78376 403678 78432
rect 344926 4120 344982 4176
rect 349710 3984 349766 4040
rect 356150 3984 356206 4040
rect 356334 3984 356390 4040
rect 398102 3984 398158 4040
rect 398286 3984 398342 4040
rect 349986 3848 350042 3904
rect 344926 3712 344982 3768
rect 339682 3168 339738 3224
rect 356150 3168 356206 3224
rect 398102 3168 398158 3224
rect 407762 77832 407818 77888
rect 407762 77424 407818 77480
rect 414662 78512 414718 78568
rect 413466 77832 413522 77888
rect 411994 77560 412050 77616
rect 410338 77288 410394 77344
rect 418158 77968 418214 78024
rect 416594 77560 416650 77616
rect 415030 77424 415086 77480
rect 414662 3984 414718 4040
rect 411994 3576 412050 3632
rect 422850 78512 422906 78568
rect 421286 77696 421342 77752
rect 432234 78512 432290 78568
rect 435362 9016 435418 9072
rect 433798 8880 433854 8936
rect 429106 5344 429162 5400
rect 427542 5072 427598 5128
rect 425978 4936 426034 4992
rect 443182 9560 443238 9616
rect 441618 9424 441674 9480
rect 440054 9288 440110 9344
rect 438490 9152 438546 9208
rect 446310 78104 446366 78160
rect 444746 8608 444802 8664
rect 449438 78240 449494 78296
rect 447874 4800 447930 4856
rect 436926 4664 436982 4720
rect 452566 78376 452622 78432
rect 451002 3848 451058 3904
rect 419722 3440 419778 3496
rect 403622 3168 403678 3224
rect 398286 3032 398342 3088
<< metal3 >>
rect 192334 700436 192340 700500
rect 192404 700498 192410 700500
rect 348785 700498 348851 700501
rect 192404 700496 348851 700498
rect 192404 700440 348790 700496
rect 348846 700440 348851 700496
rect 192404 700438 348851 700440
rect 192404 700436 192410 700438
rect 348785 700435 348851 700438
rect 109033 700362 109099 700365
rect 527173 700362 527239 700365
rect 109033 700360 527239 700362
rect 109033 700304 109038 700360
rect 109094 700304 527178 700360
rect 527234 700304 527239 700360
rect 109033 700302 527239 700304
rect 109033 700299 109099 700302
rect 527173 700299 527239 700302
rect -960 697220 480 697460
rect 104709 697234 104775 697237
rect 583520 697234 584960 697324
rect 104709 697232 584960 697234
rect 104709 697176 104714 697232
rect 104770 697176 584960 697232
rect 104709 697174 584960 697176
rect 104709 697171 104775 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 100385 644058 100451 644061
rect 583520 644058 584960 644148
rect 100385 644056 584960 644058
rect 100385 644000 100390 644056
rect 100446 644000 584960 644056
rect 100385 643998 584960 644000
rect 100385 643995 100451 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 152273 630866 152339 630869
rect 583520 630866 584960 630956
rect 152273 630864 584960 630866
rect 152273 630808 152278 630864
rect 152334 630808 584960 630864
rect 152273 630806 584960 630808
rect 152273 630803 152339 630806
rect 583520 630716 584960 630806
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 96061 591018 96127 591021
rect 583520 591018 584960 591108
rect 96061 591016 584960 591018
rect 96061 590960 96066 591016
rect 96122 590960 584960 591016
rect 96061 590958 584960 590960
rect 96061 590955 96127 590958
rect 583520 590868 584960 590958
rect -960 579852 480 580092
rect 147949 577690 148015 577693
rect 583520 577690 584960 577780
rect 147949 577688 584960 577690
rect 147949 577632 147954 577688
rect 148010 577632 584960 577688
rect 147949 577630 584960 577632
rect 147949 577627 148015 577630
rect 583520 577540 584960 577630
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 91737 537842 91803 537845
rect 583520 537842 584960 537932
rect 91737 537840 584960 537842
rect 91737 537784 91742 537840
rect 91798 537784 584960 537840
rect 91737 537782 584960 537784
rect 91737 537779 91803 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 143625 524514 143691 524517
rect 583520 524514 584960 524604
rect 143625 524512 584960 524514
rect 143625 524456 143630 524512
rect 143686 524456 584960 524512
rect 143625 524454 584960 524456
rect 143625 524451 143691 524454
rect 583520 524364 584960 524454
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 87413 484666 87479 484669
rect 583520 484666 584960 484756
rect 87413 484664 584960 484666
rect 87413 484608 87418 484664
rect 87474 484608 584960 484664
rect 87413 484606 584960 484608
rect 87413 484603 87479 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 139301 471474 139367 471477
rect 583520 471474 584960 471564
rect 139301 471472 584960 471474
rect 139301 471416 139306 471472
rect 139362 471416 584960 471472
rect 139301 471414 584960 471416
rect 139301 471411 139367 471414
rect 583520 471324 584960 471414
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 83089 298754 83155 298757
rect 583520 298754 584960 298844
rect 83089 298752 584960 298754
rect 83089 298696 83094 298752
rect 83150 298696 584960 298752
rect 83089 298694 584960 298696
rect 83089 298691 83155 298694
rect 583520 298604 584960 298694
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 118049 192674 118115 192677
rect 397453 192674 397519 192677
rect 118049 192672 397519 192674
rect 118049 192616 118054 192672
rect 118110 192616 397458 192672
rect 397514 192616 397519 192672
rect 118049 192614 397519 192616
rect 118049 192611 118115 192614
rect 397453 192611 397519 192614
rect 113633 192538 113699 192541
rect 462313 192538 462379 192541
rect 113633 192536 462379 192538
rect 113633 192480 113638 192536
rect 113694 192480 462318 192536
rect 462374 192480 462379 192536
rect 113633 192478 462379 192480
rect 113633 192475 113699 192478
rect 462313 192475 462379 192478
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 191833 186554 191899 186557
rect 189796 186552 191899 186554
rect 189796 186496 191838 186552
rect 191894 186496 191899 186552
rect 189796 186494 191899 186496
rect 191833 186491 191899 186494
rect 191925 183426 191991 183429
rect 189796 183424 191991 183426
rect 189796 183368 191930 183424
rect 191986 183368 191991 183424
rect 189796 183366 191991 183368
rect 191925 183363 191991 183366
rect 192017 180298 192083 180301
rect 189796 180296 192083 180298
rect 189796 180240 192022 180296
rect 192078 180240 192083 180296
rect 189796 180238 192083 180240
rect 192017 180235 192083 180238
rect 583520 179060 584960 179300
rect 191782 177170 191788 177172
rect 189796 177110 191788 177170
rect 191782 177108 191788 177110
rect 191852 177108 191858 177172
rect -960 175796 480 176036
rect 192109 174042 192175 174045
rect 189796 174040 192175 174042
rect 189796 173984 192114 174040
rect 192170 173984 192175 174040
rect 189796 173982 192175 173984
rect 192109 173979 192175 173982
rect 192201 170914 192267 170917
rect 189796 170912 192267 170914
rect 189796 170856 192206 170912
rect 192262 170856 192267 170912
rect 189796 170854 192267 170856
rect 192201 170851 192267 170854
rect 192293 167786 192359 167789
rect 189796 167784 192359 167786
rect 189796 167728 192298 167784
rect 192354 167728 192359 167784
rect 189796 167726 192359 167728
rect 192293 167723 192359 167726
rect 583520 165732 584960 165972
rect 190453 164658 190519 164661
rect 189796 164656 190519 164658
rect 189796 164600 190458 164656
rect 190514 164600 190519 164656
rect 189796 164598 190519 164600
rect 190453 164595 190519 164598
rect -960 162740 480 162980
rect 190545 161530 190611 161533
rect 189796 161528 190611 161530
rect 189796 161472 190550 161528
rect 190606 161472 190611 161528
rect 189796 161470 190611 161472
rect 190545 161467 190611 161470
rect 192385 158402 192451 158405
rect 189796 158400 192451 158402
rect 189796 158344 192390 158400
rect 192446 158344 192451 158400
rect 189796 158342 192451 158344
rect 192385 158339 192451 158342
rect 192477 155274 192543 155277
rect 189796 155272 192543 155274
rect 189796 155216 192482 155272
rect 192538 155216 192543 155272
rect 189796 155214 192543 155216
rect 192477 155211 192543 155214
rect 583520 152540 584960 152780
rect 190637 152146 190703 152149
rect 189796 152144 190703 152146
rect 189796 152088 190642 152144
rect 190698 152088 190703 152144
rect 189796 152086 190703 152088
rect 190637 152083 190703 152086
rect -960 149684 480 149924
rect 192569 149018 192635 149021
rect 189796 149016 192635 149018
rect 189796 148960 192574 149016
rect 192630 148960 192635 149016
rect 189796 148958 192635 148960
rect 192569 148955 192635 148958
rect 190729 145890 190795 145893
rect 189796 145888 190795 145890
rect 189796 145832 190734 145888
rect 190790 145832 190795 145888
rect 189796 145830 190795 145832
rect 190729 145827 190795 145830
rect 190821 142762 190887 142765
rect 189796 142760 190887 142762
rect 189796 142704 190826 142760
rect 190882 142704 190887 142760
rect 189796 142702 190887 142704
rect 190821 142699 190887 142702
rect 190913 139634 190979 139637
rect 189796 139632 190979 139634
rect 189796 139576 190918 139632
rect 190974 139576 190979 139632
rect 189796 139574 190979 139576
rect 190913 139571 190979 139574
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 189766 135826 189826 136476
rect 189993 135826 190059 135829
rect 189766 135824 190059 135826
rect 189766 135768 189998 135824
rect 190054 135768 190059 135824
rect 189766 135766 190059 135768
rect 189993 135763 190059 135766
rect 191005 133378 191071 133381
rect 189796 133376 191071 133378
rect 189796 133320 191010 133376
rect 191066 133320 191071 133376
rect 189796 133318 191071 133320
rect 191005 133315 191071 133318
rect 191097 130250 191163 130253
rect 189796 130248 191163 130250
rect 189796 130192 191102 130248
rect 191158 130192 191163 130248
rect 189796 130190 191163 130192
rect 191097 130187 191163 130190
rect 191230 127122 191236 127124
rect 189796 127062 191236 127122
rect 191230 127060 191236 127062
rect 191300 127060 191306 127124
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 189398 123453 189458 123964
rect 189349 123448 189458 123453
rect 189349 123392 189354 123448
rect 189410 123392 189458 123448
rect 189349 123390 189458 123392
rect 189349 123387 189415 123390
rect 189398 120325 189458 120836
rect 267733 120594 267799 120597
rect 304533 120594 304599 120597
rect 267733 120592 304599 120594
rect 267733 120536 267738 120592
rect 267794 120536 304538 120592
rect 304594 120536 304599 120592
rect 267733 120534 304599 120536
rect 267733 120531 267799 120534
rect 304533 120531 304599 120534
rect 271229 120458 271295 120461
rect 313641 120458 313707 120461
rect 271229 120456 313707 120458
rect 271229 120400 271234 120456
rect 271290 120400 313646 120456
rect 313702 120400 313707 120456
rect 271229 120398 313707 120400
rect 271229 120395 271295 120398
rect 313641 120395 313707 120398
rect 189398 120320 189507 120325
rect 189398 120264 189446 120320
rect 189502 120264 189507 120320
rect 189398 120262 189507 120264
rect 189441 120259 189507 120262
rect 274817 120322 274883 120325
rect 322749 120322 322815 120325
rect 274817 120320 322815 120322
rect 274817 120264 274822 120320
rect 274878 120264 322754 120320
rect 322810 120264 322815 120320
rect 274817 120262 322815 120264
rect 274817 120259 274883 120262
rect 322749 120259 322815 120262
rect 264145 120186 264211 120189
rect 331857 120186 331923 120189
rect 264145 120184 331923 120186
rect 264145 120128 264150 120184
rect 264206 120128 331862 120184
rect 331918 120128 331923 120184
rect 264145 120126 331923 120128
rect 264145 120123 264211 120126
rect 331857 120123 331923 120126
rect 191189 117738 191255 117741
rect 189796 117736 191255 117738
rect 189796 117680 191194 117736
rect 191250 117680 191255 117736
rect 189796 117678 191255 117680
rect 191189 117675 191255 117678
rect 335854 117404 335860 117468
rect 335924 117404 335930 117468
rect 336038 116452 336044 116516
rect 336108 116452 336114 116516
rect 339769 115562 339835 115565
rect 336260 115560 339835 115562
rect 336260 115504 339774 115560
rect 339830 115504 339835 115560
rect 336260 115502 339835 115504
rect 339769 115499 339835 115502
rect 190494 114610 190500 114612
rect 189796 114550 190500 114610
rect 190494 114548 190500 114550
rect 190564 114548 190570 114612
rect 338113 114610 338179 114613
rect 336260 114608 338179 114610
rect 336260 114552 338118 114608
rect 338174 114552 338179 114608
rect 336260 114550 338179 114552
rect 338113 114547 338179 114550
rect 339493 113658 339559 113661
rect 336260 113656 339559 113658
rect 336260 113600 339498 113656
rect 339554 113600 339559 113656
rect 336260 113598 339559 113600
rect 339493 113595 339559 113598
rect 337469 112706 337535 112709
rect 336260 112704 337535 112706
rect 336260 112648 337474 112704
rect 337530 112648 337535 112704
rect 583520 112692 584960 112932
rect 336260 112646 337535 112648
rect 337469 112643 337535 112646
rect 338982 111754 338988 111756
rect 336260 111694 338988 111754
rect 338982 111692 338988 111694
rect 339052 111692 339058 111756
rect 189582 110941 189642 111452
rect 189533 110936 189642 110941
rect 189533 110880 189538 110936
rect 189594 110880 189642 110936
rect 189533 110878 189642 110880
rect 189533 110875 189599 110878
rect 336774 110802 336780 110804
rect -960 110516 480 110756
rect 336260 110742 336780 110802
rect 336774 110740 336780 110742
rect 336844 110740 336850 110804
rect 338614 109850 338620 109852
rect 336260 109790 338620 109850
rect 338614 109788 338620 109790
rect 338684 109788 338690 109852
rect 336046 108357 336106 108868
rect 192661 108354 192727 108357
rect 189796 108352 192727 108354
rect 189796 108296 192666 108352
rect 192722 108296 192727 108352
rect 189796 108294 192727 108296
rect 192661 108291 192727 108294
rect 335997 108352 336106 108357
rect 335997 108296 336002 108352
rect 336058 108296 336106 108352
rect 335997 108294 336106 108296
rect 335997 108291 336063 108294
rect 336222 107884 336228 107948
rect 336292 107884 336298 107948
rect 398097 107810 398163 107813
rect 398097 107808 400108 107810
rect 398097 107752 398102 107808
rect 398158 107752 400108 107808
rect 398097 107750 400108 107752
rect 398097 107747 398163 107750
rect 336825 106994 336891 106997
rect 336260 106992 336891 106994
rect 336260 106936 336830 106992
rect 336886 106936 336891 106992
rect 336260 106934 336891 106936
rect 336825 106931 336891 106934
rect 338430 106042 338436 106044
rect 336260 105982 338436 106042
rect 338430 105980 338436 105982
rect 338500 105980 338506 106044
rect 191281 105226 191347 105229
rect 189796 105224 191347 105226
rect 189796 105168 191286 105224
rect 191342 105168 191347 105224
rect 189796 105166 191347 105168
rect 191281 105163 191347 105166
rect 336733 105090 336799 105093
rect 336260 105088 336799 105090
rect 336260 105032 336738 105088
rect 336794 105032 336799 105088
rect 336260 105030 336799 105032
rect 336733 105027 336799 105030
rect 338297 104138 338363 104141
rect 336260 104136 338363 104138
rect 336260 104080 338302 104136
rect 338358 104080 338363 104136
rect 336260 104078 338363 104080
rect 338297 104075 338363 104078
rect 336917 103186 336983 103189
rect 336260 103184 336983 103186
rect 336260 103128 336922 103184
rect 336978 103128 336983 103184
rect 336260 103126 336983 103128
rect 336917 103123 336983 103126
rect 338205 102234 338271 102237
rect 336260 102232 338271 102234
rect 336260 102176 338210 102232
rect 338266 102176 338271 102232
rect 336260 102174 338271 102176
rect 338205 102171 338271 102174
rect 189582 101557 189642 102068
rect 189582 101552 189691 101557
rect 189582 101496 189630 101552
rect 189686 101496 189691 101552
rect 189582 101494 189691 101496
rect 189625 101491 189691 101494
rect 337377 101282 337443 101285
rect 336260 101280 337443 101282
rect 336260 101224 337382 101280
rect 337438 101224 337443 101280
rect 336260 101222 337443 101224
rect 337377 101219 337443 101222
rect 339585 100330 339651 100333
rect 336260 100328 339651 100330
rect 336260 100272 339590 100328
rect 339646 100272 339651 100328
rect 336260 100270 339651 100272
rect 339585 100267 339651 100270
rect 583520 99364 584960 99604
rect 189390 98908 189396 98972
rect 189460 98908 189466 98972
rect 336230 98698 336290 99348
rect 336406 98698 336412 98700
rect 336230 98638 336412 98698
rect 336406 98636 336412 98638
rect 336476 98636 336482 98700
rect 338798 98426 338804 98428
rect 336260 98366 338804 98426
rect 338798 98364 338804 98366
rect 338868 98364 338874 98428
rect -960 97460 480 97700
rect 336046 96933 336106 97444
rect 336046 96928 336155 96933
rect 336046 96872 336094 96928
rect 336150 96872 336155 96928
rect 336046 96870 336155 96872
rect 336089 96867 336155 96870
rect 338849 96522 338915 96525
rect 336260 96520 338915 96522
rect 336260 96464 338854 96520
rect 338910 96464 338915 96520
rect 336260 96462 338915 96464
rect 338849 96459 338915 96462
rect 189766 95298 189826 95812
rect 337009 95570 337075 95573
rect 336260 95568 337075 95570
rect 336260 95512 337014 95568
rect 337070 95512 337075 95568
rect 336260 95510 337075 95512
rect 337009 95507 337075 95510
rect 189901 95298 189967 95301
rect 189766 95296 189967 95298
rect 189766 95240 189906 95296
rect 189962 95240 189967 95296
rect 189766 95238 189967 95240
rect 189901 95235 189967 95238
rect 338481 94618 338547 94621
rect 336260 94616 338547 94618
rect 336260 94560 338486 94616
rect 338542 94560 338547 94616
rect 336260 94558 338547 94560
rect 338481 94555 338547 94558
rect 337101 93666 337167 93669
rect 336260 93664 337167 93666
rect 336260 93608 337106 93664
rect 337162 93608 337167 93664
rect 336260 93606 337167 93608
rect 337101 93603 337167 93606
rect 190862 92714 190868 92716
rect 189796 92654 190868 92714
rect 190862 92652 190868 92654
rect 190932 92652 190938 92716
rect 338389 92714 338455 92717
rect 336260 92712 338455 92714
rect 336260 92656 338394 92712
rect 338450 92656 338455 92712
rect 336260 92654 338455 92656
rect 338389 92651 338455 92654
rect 337193 91762 337259 91765
rect 336260 91760 337259 91762
rect 336260 91704 337198 91760
rect 337254 91704 337259 91760
rect 336260 91702 337259 91704
rect 337193 91699 337259 91702
rect 338573 90810 338639 90813
rect 336260 90808 338639 90810
rect 336260 90752 338578 90808
rect 338634 90752 338639 90808
rect 336260 90750 338639 90752
rect 338573 90747 338639 90750
rect 336230 89589 336290 89828
rect 336230 89584 336339 89589
rect 189766 88909 189826 89556
rect 336230 89528 336278 89584
rect 336334 89528 336339 89584
rect 336230 89526 336339 89528
rect 336273 89523 336339 89526
rect 189766 88904 189875 88909
rect 189766 88848 189814 88904
rect 189870 88848 189875 88904
rect 189766 88846 189875 88848
rect 189809 88843 189875 88846
rect 336230 88365 336290 88876
rect 336181 88360 336290 88365
rect 336181 88304 336186 88360
rect 336242 88304 336290 88360
rect 336181 88302 336290 88304
rect 336181 88299 336247 88302
rect 336230 87274 336290 87924
rect 336365 87274 336431 87277
rect 336230 87272 336431 87274
rect 336230 87216 336370 87272
rect 336426 87216 336431 87272
rect 336230 87214 336431 87216
rect 336365 87211 336431 87214
rect 338757 87002 338823 87005
rect 336260 87000 338823 87002
rect 336260 86944 338762 87000
rect 338818 86944 338823 87000
rect 336260 86942 338823 86944
rect 338757 86939 338823 86942
rect 192334 86458 192340 86460
rect 189796 86398 192340 86458
rect 192334 86396 192340 86398
rect 192404 86396 192410 86460
rect 337285 86050 337351 86053
rect 336260 86048 337351 86050
rect 336260 85992 337290 86048
rect 337346 85992 337351 86048
rect 583520 86036 584960 86276
rect 336260 85990 337351 85992
rect 337285 85987 337351 85990
rect 338941 85098 339007 85101
rect 336260 85096 339007 85098
rect 336260 85040 338946 85096
rect 339002 85040 339007 85096
rect 336260 85038 339007 85040
rect 338941 85035 339007 85038
rect -960 84540 480 84780
rect 339677 84146 339743 84149
rect 336260 84144 339743 84146
rect 336260 84088 339682 84144
rect 339738 84088 339743 84144
rect 336260 84086 339743 84088
rect 339677 84083 339743 84086
rect 191966 83330 191972 83332
rect 189796 83270 191972 83330
rect 191966 83268 191972 83270
rect 192036 83268 192042 83332
rect 338297 83194 338363 83197
rect 336260 83192 338363 83194
rect 336260 83136 338302 83192
rect 338358 83136 338363 83192
rect 336260 83134 338363 83136
rect 338297 83131 338363 83134
rect 336230 81562 336290 82212
rect 336549 81562 336615 81565
rect 336230 81560 336615 81562
rect 336230 81504 336554 81560
rect 336610 81504 336615 81560
rect 336230 81502 336615 81504
rect 336549 81499 336615 81502
rect 335670 81228 335676 81292
rect 335740 81228 335746 81292
rect 338665 81154 338731 81157
rect 338070 81152 338731 81154
rect 338070 81096 338670 81152
rect 338726 81096 338731 81152
rect 338070 81094 338731 81096
rect 193857 80746 193923 80749
rect 338070 80746 338130 81094
rect 338665 81091 338731 81094
rect 193857 80744 338130 80746
rect 193857 80688 193862 80744
rect 193918 80688 338130 80744
rect 193857 80686 338130 80688
rect 193857 80683 193923 80686
rect 189717 80610 189783 80613
rect 335670 80610 335676 80612
rect 189717 80608 335676 80610
rect 189717 80552 189722 80608
rect 189778 80552 335676 80608
rect 189717 80550 335676 80552
rect 189717 80547 189783 80550
rect 335670 80548 335676 80550
rect 335740 80548 335746 80612
rect 336641 80066 336707 80069
rect 315990 80064 336707 80066
rect 315990 80008 336646 80064
rect 336702 80008 336707 80064
rect 315990 80006 336707 80008
rect 246389 79658 246455 79661
rect 315990 79658 316050 80006
rect 336641 80003 336707 80006
rect 246389 79656 316050 79658
rect 246389 79600 246394 79656
rect 246450 79600 316050 79656
rect 246389 79598 316050 79600
rect 246389 79595 246455 79598
rect 207381 79522 207447 79525
rect 339769 79522 339835 79525
rect 207381 79520 339835 79522
rect 207381 79464 207386 79520
rect 207442 79464 339774 79520
rect 339830 79464 339835 79520
rect 207381 79462 339835 79464
rect 207381 79459 207447 79462
rect 339769 79459 339835 79462
rect 168373 79386 168439 79389
rect 338297 79386 338363 79389
rect 168373 79384 338363 79386
rect 168373 79328 168378 79384
rect 168434 79328 338302 79384
rect 338358 79328 338363 79384
rect 168373 79326 338363 79328
rect 168373 79323 168439 79326
rect 338297 79323 338363 79326
rect 105721 78570 105787 78573
rect 180241 78570 180307 78573
rect 105721 78568 180307 78570
rect 105721 78512 105726 78568
rect 105782 78512 180246 78568
rect 180302 78512 180307 78568
rect 105721 78510 180307 78512
rect 105721 78507 105787 78510
rect 180241 78507 180307 78510
rect 324262 78508 324268 78572
rect 324332 78570 324338 78572
rect 324957 78570 325023 78573
rect 324332 78568 325023 78570
rect 324332 78512 324962 78568
rect 325018 78512 325023 78568
rect 324332 78510 325023 78512
rect 324332 78508 324338 78510
rect 324957 78507 325023 78510
rect 414657 78570 414723 78573
rect 422845 78570 422911 78573
rect 414657 78568 422911 78570
rect 414657 78512 414662 78568
rect 414718 78512 422850 78568
rect 422906 78512 422911 78568
rect 414657 78510 422911 78512
rect 414657 78507 414723 78510
rect 422845 78507 422911 78510
rect 431902 78508 431908 78572
rect 431972 78570 431978 78572
rect 432229 78570 432295 78573
rect 431972 78568 432295 78570
rect 431972 78512 432234 78568
rect 432290 78512 432295 78568
rect 431972 78510 432295 78512
rect 431972 78508 431978 78510
rect 432229 78507 432295 78510
rect 178677 78434 178743 78437
rect 171182 78432 178743 78434
rect 171182 78376 178682 78432
rect 178738 78376 178743 78432
rect 171182 78374 178743 78376
rect 91553 78298 91619 78301
rect 124121 78298 124187 78301
rect 91553 78296 124187 78298
rect 91553 78240 91558 78296
rect 91614 78240 124126 78296
rect 124182 78240 124187 78296
rect 91553 78238 124187 78240
rect 91553 78235 91619 78238
rect 124121 78235 124187 78238
rect 116117 78162 116183 78165
rect 118693 78162 118759 78165
rect 116117 78160 118759 78162
rect 116117 78104 116122 78160
rect 116178 78104 118698 78160
rect 118754 78104 118759 78160
rect 116117 78102 118759 78104
rect 116117 78099 116183 78102
rect 118693 78099 118759 78102
rect 162894 78100 162900 78164
rect 162964 78162 162970 78164
rect 163037 78162 163103 78165
rect 162964 78160 163103 78162
rect 162964 78104 163042 78160
rect 163098 78104 163103 78160
rect 162964 78102 163103 78104
rect 162964 78100 162970 78102
rect 163037 78099 163103 78102
rect 4061 78026 4127 78029
rect 84837 78026 84903 78029
rect 4061 78024 84903 78026
rect 4061 77968 4066 78024
rect 4122 77968 84842 78024
rect 84898 77968 84903 78024
rect 4061 77966 84903 77968
rect 4061 77963 4127 77966
rect 84837 77963 84903 77966
rect 102225 78026 102291 78029
rect 171182 78026 171242 78374
rect 178677 78371 178743 78374
rect 179229 78434 179295 78437
rect 306925 78434 306991 78437
rect 179229 78432 306991 78434
rect 179229 78376 179234 78432
rect 179290 78376 306930 78432
rect 306986 78376 306991 78432
rect 179229 78374 306991 78376
rect 179229 78371 179295 78374
rect 306925 78371 306991 78374
rect 403617 78434 403683 78437
rect 452561 78434 452627 78437
rect 403617 78432 452627 78434
rect 403617 78376 403622 78432
rect 403678 78376 452566 78432
rect 452622 78376 452627 78432
rect 403617 78374 452627 78376
rect 403617 78371 403683 78374
rect 452561 78371 452627 78374
rect 180057 78298 180123 78301
rect 315941 78298 316007 78301
rect 180057 78296 316007 78298
rect 180057 78240 180062 78296
rect 180118 78240 315946 78296
rect 316002 78240 316007 78296
rect 180057 78238 316007 78240
rect 180057 78235 180123 78238
rect 315941 78235 316007 78238
rect 335077 78298 335143 78301
rect 449433 78298 449499 78301
rect 335077 78296 449499 78298
rect 335077 78240 335082 78296
rect 335138 78240 449438 78296
rect 449494 78240 449499 78296
rect 335077 78238 449499 78240
rect 335077 78235 335143 78238
rect 449433 78235 449499 78238
rect 178953 78162 179019 78165
rect 320449 78162 320515 78165
rect 178953 78160 320515 78162
rect 178953 78104 178958 78160
rect 179014 78104 320454 78160
rect 320510 78104 320515 78160
rect 178953 78102 320515 78104
rect 178953 78099 179019 78102
rect 320449 78099 320515 78102
rect 327993 78162 328059 78165
rect 446305 78162 446371 78165
rect 327993 78160 446371 78162
rect 327993 78104 327998 78160
rect 328054 78104 446310 78160
rect 446366 78104 446371 78160
rect 327993 78102 446371 78104
rect 327993 78099 328059 78102
rect 446305 78099 446371 78102
rect 177113 78026 177179 78029
rect 102225 78024 171242 78026
rect 102225 77968 102230 78024
rect 102286 77968 171242 78024
rect 102225 77966 171242 77968
rect 174310 78024 177179 78026
rect 174310 77968 177118 78024
rect 177174 77968 177179 78024
rect 174310 77966 177179 77968
rect 102225 77963 102291 77966
rect 5257 77890 5323 77893
rect 86401 77890 86467 77893
rect 5257 77888 86467 77890
rect 5257 77832 5262 77888
rect 5318 77832 86406 77888
rect 86462 77832 86467 77888
rect 5257 77830 86467 77832
rect 5257 77827 5323 77830
rect 86401 77827 86467 77830
rect 98637 77890 98703 77893
rect 144913 77890 144979 77893
rect 98637 77888 144979 77890
rect 98637 77832 98642 77888
rect 98698 77832 144918 77888
rect 144974 77832 144979 77888
rect 98637 77830 144979 77832
rect 98637 77827 98703 77830
rect 144913 77827 144979 77830
rect 145046 77828 145052 77892
rect 145116 77890 145122 77892
rect 145833 77890 145899 77893
rect 145116 77888 145899 77890
rect 145116 77832 145838 77888
rect 145894 77832 145899 77888
rect 145116 77830 145899 77832
rect 145116 77828 145122 77830
rect 145833 77827 145899 77830
rect 146017 77890 146083 77893
rect 174310 77890 174370 77966
rect 177113 77963 177179 77966
rect 222745 78026 222811 78029
rect 418153 78026 418219 78029
rect 222745 78024 418219 78026
rect 222745 77968 222750 78024
rect 222806 77968 418158 78024
rect 418214 77968 418219 78024
rect 222745 77966 418219 77968
rect 222745 77963 222811 77966
rect 418153 77963 418219 77966
rect 146017 77888 174370 77890
rect 146017 77832 146022 77888
rect 146078 77832 174370 77888
rect 146017 77830 174370 77832
rect 146017 77827 146083 77830
rect 175222 77828 175228 77892
rect 175292 77890 175298 77892
rect 175549 77890 175615 77893
rect 175292 77888 175615 77890
rect 175292 77832 175554 77888
rect 175610 77832 175615 77888
rect 175292 77830 175615 77832
rect 175292 77828 175298 77830
rect 175549 77827 175615 77830
rect 215661 77890 215727 77893
rect 407757 77890 407823 77893
rect 215661 77888 407823 77890
rect 215661 77832 215666 77888
rect 215722 77832 407762 77888
rect 407818 77832 407823 77888
rect 215661 77830 407823 77832
rect 215661 77827 215727 77830
rect 407757 77827 407823 77830
rect 410374 77828 410380 77892
rect 410444 77890 410450 77892
rect 413461 77890 413527 77893
rect 410444 77888 413527 77890
rect 410444 77832 413466 77888
rect 413522 77832 413527 77888
rect 410444 77830 413527 77832
rect 410444 77828 410450 77830
rect 413461 77827 413527 77830
rect 112805 77754 112871 77757
rect 183369 77754 183435 77757
rect 112805 77752 183435 77754
rect 112805 77696 112810 77752
rect 112866 77696 183374 77752
rect 183430 77696 183435 77752
rect 112805 77694 183435 77696
rect 112805 77691 112871 77694
rect 183369 77691 183435 77694
rect 300117 77754 300183 77757
rect 421281 77754 421347 77757
rect 300117 77752 421347 77754
rect 300117 77696 300122 77752
rect 300178 77696 421286 77752
rect 421342 77696 421347 77752
rect 300117 77694 421347 77696
rect 300117 77691 300183 77694
rect 421281 77691 421347 77694
rect 116117 77618 116183 77621
rect 84150 77558 93870 77618
rect 41873 77482 41939 77485
rect 84150 77482 84210 77558
rect 93810 77482 93870 77558
rect 103470 77616 116183 77618
rect 103470 77560 116122 77616
rect 116178 77560 116183 77616
rect 103470 77558 116183 77560
rect 103470 77482 103530 77558
rect 116117 77555 116183 77558
rect 116393 77618 116459 77621
rect 184933 77618 184999 77621
rect 116393 77616 184999 77618
rect 116393 77560 116398 77616
rect 116454 77560 184938 77616
rect 184994 77560 184999 77616
rect 116393 77558 184999 77560
rect 116393 77555 116459 77558
rect 184933 77555 184999 77558
rect 210969 77618 211035 77621
rect 336733 77618 336799 77621
rect 210969 77616 336799 77618
rect 210969 77560 210974 77616
rect 211030 77560 336738 77616
rect 336794 77560 336799 77616
rect 210969 77558 336799 77560
rect 210969 77555 211035 77558
rect 336733 77555 336799 77558
rect 411989 77618 412055 77621
rect 416589 77618 416655 77621
rect 411989 77616 416655 77618
rect 411989 77560 411994 77616
rect 412050 77560 416594 77616
rect 416650 77560 416655 77616
rect 411989 77558 416655 77560
rect 411989 77555 412055 77558
rect 416589 77555 416655 77558
rect 117221 77482 117287 77485
rect 41873 77480 84210 77482
rect 41873 77424 41878 77480
rect 41934 77424 84210 77480
rect 41873 77422 84210 77424
rect 88934 77422 91386 77482
rect 93810 77422 103530 77482
rect 114510 77480 117287 77482
rect 114510 77424 117226 77480
rect 117282 77424 117287 77480
rect 114510 77422 117287 77424
rect 41873 77419 41939 77422
rect 18229 77346 18295 77349
rect 88934 77346 88994 77422
rect 18229 77344 88994 77346
rect 18229 77288 18234 77344
rect 18290 77288 88994 77344
rect 18229 77286 88994 77288
rect 91093 77348 91159 77349
rect 91093 77344 91140 77348
rect 91204 77346 91210 77348
rect 91326 77346 91386 77422
rect 114510 77346 114570 77422
rect 117221 77419 117287 77422
rect 119889 77482 119955 77485
rect 186497 77482 186563 77485
rect 119889 77480 186563 77482
rect 119889 77424 119894 77480
rect 119950 77424 186502 77480
rect 186558 77424 186563 77480
rect 119889 77422 186563 77424
rect 119889 77419 119955 77422
rect 186497 77419 186563 77422
rect 407757 77482 407823 77485
rect 415025 77482 415091 77485
rect 407757 77480 415091 77482
rect 407757 77424 407762 77480
rect 407818 77424 415030 77480
rect 415086 77424 415091 77480
rect 407757 77422 415091 77424
rect 407757 77419 407823 77422
rect 415025 77419 415091 77422
rect 91093 77288 91098 77344
rect 18229 77283 18295 77286
rect 91093 77284 91140 77288
rect 91204 77286 91250 77346
rect 91326 77286 114570 77346
rect 114645 77346 114711 77349
rect 114870 77346 114876 77348
rect 114645 77344 114876 77346
rect 114645 77288 114650 77344
rect 114706 77288 114876 77344
rect 114645 77286 114876 77288
rect 91204 77284 91210 77286
rect 91093 77283 91159 77284
rect 114645 77283 114711 77286
rect 114870 77284 114876 77286
rect 114940 77284 114946 77348
rect 123477 77346 123543 77349
rect 188061 77346 188127 77349
rect 123477 77344 188127 77346
rect 123477 77288 123482 77344
rect 123538 77288 188066 77344
rect 188122 77288 188127 77344
rect 123477 77286 188127 77288
rect 123477 77283 123543 77286
rect 188061 77283 188127 77286
rect 409086 77284 409092 77348
rect 409156 77346 409162 77348
rect 410333 77346 410399 77349
rect 409156 77344 410399 77346
rect 409156 77288 410338 77344
rect 410394 77288 410399 77344
rect 409156 77286 410399 77288
rect 409156 77284 409162 77286
rect 410333 77283 410399 77286
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 218053 22674 218119 22677
rect 337377 22674 337443 22677
rect 218053 22672 337443 22674
rect 218053 22616 218058 22672
rect 218114 22616 337382 22672
rect 337438 22616 337443 22672
rect 218053 22614 337443 22616
rect 218053 22611 218119 22614
rect 337377 22611 337443 22614
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 67909 13018 67975 13021
rect 189993 13018 190059 13021
rect 67909 13016 190059 13018
rect 67909 12960 67914 13016
rect 67970 12960 189998 13016
rect 190054 12960 190059 13016
rect 67909 12958 190059 12960
rect 67909 12955 67975 12958
rect 189993 12955 190059 12958
rect 74993 12338 75059 12341
rect 190821 12338 190887 12341
rect 74993 12336 190887 12338
rect 74993 12280 74998 12336
rect 75054 12280 190826 12336
rect 190882 12280 190887 12336
rect 74993 12278 190887 12280
rect 74993 12275 75059 12278
rect 190821 12275 190887 12278
rect 71497 12202 71563 12205
rect 190913 12202 190979 12205
rect 71497 12200 190979 12202
rect 71497 12144 71502 12200
rect 71558 12144 190918 12200
rect 190974 12144 190979 12200
rect 71497 12142 190979 12144
rect 71497 12139 71563 12142
rect 190913 12139 190979 12142
rect 64321 12066 64387 12069
rect 191005 12066 191071 12069
rect 64321 12064 191071 12066
rect 64321 12008 64326 12064
rect 64382 12008 191010 12064
rect 191066 12008 191071 12064
rect 64321 12006 191071 12008
rect 64321 12003 64387 12006
rect 191005 12003 191071 12006
rect 60825 11930 60891 11933
rect 191097 11930 191163 11933
rect 60825 11928 191163 11930
rect 60825 11872 60830 11928
rect 60886 11872 191102 11928
rect 191158 11872 191163 11928
rect 60825 11870 191163 11872
rect 60825 11867 60891 11870
rect 191097 11867 191163 11870
rect 53741 11794 53807 11797
rect 189349 11794 189415 11797
rect 53741 11792 189415 11794
rect 53741 11736 53746 11792
rect 53802 11736 189354 11792
rect 189410 11736 189415 11792
rect 53741 11734 189415 11736
rect 53741 11731 53807 11734
rect 189349 11731 189415 11734
rect 50153 11658 50219 11661
rect 189441 11658 189507 11661
rect 50153 11656 189507 11658
rect 50153 11600 50158 11656
rect 50214 11600 189446 11656
rect 189502 11600 189507 11656
rect 50153 11598 189507 11600
rect 50153 11595 50219 11598
rect 189441 11595 189507 11598
rect 78489 11522 78555 11525
rect 190729 11522 190795 11525
rect 78489 11520 190795 11522
rect 78489 11464 78494 11520
rect 78550 11464 190734 11520
rect 190790 11464 190795 11520
rect 78489 11462 190795 11464
rect 78489 11459 78555 11462
rect 190729 11459 190795 11462
rect 46657 11250 46723 11253
rect 78581 11250 78647 11253
rect 46657 11248 78647 11250
rect 46657 11192 46662 11248
rect 46718 11192 78586 11248
rect 78642 11192 78647 11248
rect 46657 11190 78647 11192
rect 46657 11187 46723 11190
rect 78581 11187 78647 11190
rect 32397 11114 32463 11117
rect 75821 11114 75887 11117
rect 32397 11112 75887 11114
rect 32397 11056 32402 11112
rect 32458 11056 75826 11112
rect 75882 11056 75887 11112
rect 32397 11054 75887 11056
rect 32397 11051 32463 11054
rect 75821 11051 75887 11054
rect 84469 10978 84535 10981
rect 170949 10978 171015 10981
rect 84469 10976 171015 10978
rect 84469 10920 84474 10976
rect 84530 10920 170954 10976
rect 171010 10920 171015 10976
rect 84469 10918 171015 10920
rect 84469 10915 84535 10918
rect 170949 10915 171015 10918
rect 80881 10842 80947 10845
rect 169385 10842 169451 10845
rect 80881 10840 169451 10842
rect 80881 10784 80886 10840
rect 80942 10784 169390 10840
rect 169446 10784 169451 10840
rect 80881 10782 169451 10784
rect 80881 10779 80947 10782
rect 169385 10779 169451 10782
rect 45461 10706 45527 10709
rect 153745 10706 153811 10709
rect 45461 10704 153811 10706
rect 45461 10648 45466 10704
rect 45522 10648 153750 10704
rect 153806 10648 153811 10704
rect 45461 10646 153811 10648
rect 45461 10643 45527 10646
rect 153745 10643 153811 10646
rect 38377 10570 38443 10573
rect 150617 10570 150683 10573
rect 38377 10568 150683 10570
rect 38377 10512 38382 10568
rect 38438 10512 150622 10568
rect 150678 10512 150683 10568
rect 38377 10510 150683 10512
rect 38377 10507 38443 10510
rect 150617 10507 150683 10510
rect 260649 10570 260715 10573
rect 336825 10570 336891 10573
rect 260649 10568 336891 10570
rect 260649 10512 260654 10568
rect 260710 10512 336830 10568
rect 336886 10512 336891 10568
rect 260649 10510 336891 10512
rect 260649 10507 260715 10510
rect 336825 10507 336891 10510
rect 34789 10434 34855 10437
rect 149053 10434 149119 10437
rect 34789 10432 149119 10434
rect 34789 10376 34794 10432
rect 34850 10376 149058 10432
rect 149114 10376 149119 10432
rect 34789 10374 149119 10376
rect 34789 10371 34855 10374
rect 149053 10371 149119 10374
rect 164877 10434 164943 10437
rect 338614 10434 338620 10436
rect 164877 10432 338620 10434
rect 164877 10376 164882 10432
rect 164938 10376 338620 10432
rect 164877 10374 338620 10376
rect 164877 10371 164943 10374
rect 338614 10372 338620 10374
rect 338684 10372 338690 10436
rect 31293 10298 31359 10301
rect 147489 10298 147555 10301
rect 31293 10296 147555 10298
rect 31293 10240 31298 10296
rect 31354 10240 147494 10296
rect 147550 10240 147555 10296
rect 31293 10238 147555 10240
rect 31293 10235 31359 10238
rect 147489 10235 147555 10238
rect 158897 10298 158963 10301
rect 338798 10298 338804 10300
rect 158897 10296 338804 10298
rect 158897 10240 158902 10296
rect 158958 10240 338804 10296
rect 158897 10238 338804 10240
rect 158897 10235 158963 10238
rect 338798 10236 338804 10238
rect 338868 10236 338874 10300
rect 87965 10162 88031 10165
rect 172513 10162 172579 10165
rect 87965 10160 172579 10162
rect 87965 10104 87970 10160
rect 88026 10104 172518 10160
rect 172574 10104 172579 10160
rect 87965 10102 172579 10104
rect 87965 10099 88031 10102
rect 172513 10099 172579 10102
rect 23013 9754 23079 9757
rect 88241 9754 88307 9757
rect 23013 9752 88307 9754
rect 23013 9696 23018 9752
rect 23074 9696 88246 9752
rect 88302 9696 88307 9752
rect 23013 9694 88307 9696
rect 23013 9691 23079 9694
rect 88241 9691 88307 9694
rect 97809 9618 97875 9621
rect 127157 9618 127223 9621
rect 97809 9616 127223 9618
rect 97809 9560 97814 9616
rect 97870 9560 127162 9616
rect 127218 9560 127223 9616
rect 97809 9558 127223 9560
rect 97809 9555 97875 9558
rect 127157 9555 127223 9558
rect 320909 9618 320975 9621
rect 443177 9618 443243 9621
rect 320909 9616 443243 9618
rect 320909 9560 320914 9616
rect 320970 9560 443182 9616
rect 443238 9560 443243 9616
rect 320909 9558 443243 9560
rect 320909 9555 320975 9558
rect 443177 9555 443243 9558
rect 93945 9482 94011 9485
rect 125593 9482 125659 9485
rect 93945 9480 125659 9482
rect 93945 9424 93950 9480
rect 94006 9424 125598 9480
rect 125654 9424 125659 9480
rect 93945 9422 125659 9424
rect 93945 9419 94011 9422
rect 125593 9419 125659 9422
rect 317229 9482 317295 9485
rect 441613 9482 441679 9485
rect 317229 9480 441679 9482
rect 317229 9424 317234 9480
rect 317290 9424 441618 9480
rect 441674 9424 441679 9480
rect 317229 9422 441679 9424
rect 317229 9419 317295 9422
rect 441613 9419 441679 9422
rect 90357 9346 90423 9349
rect 124029 9346 124095 9349
rect 90357 9344 124095 9346
rect 90357 9288 90362 9344
rect 90418 9288 124034 9344
rect 124090 9288 124095 9344
rect 90357 9286 124095 9288
rect 90357 9283 90423 9286
rect 124029 9283 124095 9286
rect 313825 9346 313891 9349
rect 440049 9346 440115 9349
rect 313825 9344 440115 9346
rect 313825 9288 313830 9344
rect 313886 9288 440054 9344
rect 440110 9288 440115 9344
rect 313825 9286 440115 9288
rect 313825 9283 313891 9286
rect 440049 9283 440115 9286
rect 44265 9210 44331 9213
rect 103697 9210 103763 9213
rect 44265 9208 103763 9210
rect 44265 9152 44270 9208
rect 44326 9152 103702 9208
rect 103758 9152 103763 9208
rect 44265 9150 103763 9152
rect 44265 9147 44331 9150
rect 103697 9147 103763 9150
rect 310237 9210 310303 9213
rect 438485 9210 438551 9213
rect 310237 9208 438551 9210
rect 310237 9152 310242 9208
rect 310298 9152 438490 9208
rect 438546 9152 438551 9208
rect 310237 9150 438551 9152
rect 310237 9147 310303 9150
rect 438485 9147 438551 9150
rect 77385 9074 77451 9077
rect 167821 9074 167887 9077
rect 77385 9072 167887 9074
rect 77385 9016 77390 9072
rect 77446 9016 167826 9072
rect 167882 9016 167887 9072
rect 77385 9014 167887 9016
rect 77385 9011 77451 9014
rect 167821 9011 167887 9014
rect 229829 9074 229895 9077
rect 300117 9074 300183 9077
rect 229829 9072 300183 9074
rect 229829 9016 229834 9072
rect 229890 9016 300122 9072
rect 300178 9016 300183 9072
rect 229829 9014 300183 9016
rect 229829 9011 229895 9014
rect 300117 9011 300183 9014
rect 303153 9074 303219 9077
rect 435357 9074 435423 9077
rect 303153 9072 435423 9074
rect 303153 9016 303158 9072
rect 303214 9016 435362 9072
rect 435418 9016 435423 9072
rect 303153 9014 435423 9016
rect 303153 9011 303219 9014
rect 435357 9011 435423 9014
rect 70301 8938 70367 8941
rect 164693 8938 164759 8941
rect 70301 8936 164759 8938
rect 70301 8880 70306 8936
rect 70362 8880 164698 8936
rect 164754 8880 164759 8936
rect 70301 8878 164759 8880
rect 70301 8875 70367 8878
rect 164693 8875 164759 8878
rect 299657 8938 299723 8941
rect 433793 8938 433859 8941
rect 299657 8936 433859 8938
rect 299657 8880 299662 8936
rect 299718 8880 433798 8936
rect 433854 8880 433859 8936
rect 299657 8878 433859 8880
rect 299657 8875 299723 8878
rect 433793 8875 433859 8878
rect 101029 8802 101095 8805
rect 128721 8802 128787 8805
rect 101029 8800 128787 8802
rect 101029 8744 101034 8800
rect 101090 8744 128726 8800
rect 128782 8744 128787 8800
rect 101029 8742 128787 8744
rect 101029 8739 101095 8742
rect 128721 8739 128787 8742
rect 292573 8802 292639 8805
rect 325601 8802 325667 8805
rect 292573 8800 325667 8802
rect 292573 8744 292578 8800
rect 292634 8744 325606 8800
rect 325662 8744 325667 8800
rect 292573 8742 325667 8744
rect 292573 8739 292639 8742
rect 325601 8739 325667 8742
rect 63217 8666 63283 8669
rect 97901 8666 97967 8669
rect 63217 8664 97967 8666
rect 63217 8608 63222 8664
rect 63278 8608 97906 8664
rect 97962 8608 97967 8664
rect 63217 8606 97967 8608
rect 63217 8603 63283 8606
rect 97901 8603 97967 8606
rect 278313 8666 278379 8669
rect 320725 8666 320791 8669
rect 278313 8664 320791 8666
rect 278313 8608 278318 8664
rect 278374 8608 320730 8664
rect 320786 8608 320791 8664
rect 278313 8606 320791 8608
rect 278313 8603 278379 8606
rect 320725 8603 320791 8606
rect 324405 8666 324471 8669
rect 444741 8666 444807 8669
rect 324405 8664 444807 8666
rect 324405 8608 324410 8664
rect 324466 8608 444746 8664
rect 444802 8608 444807 8664
rect 324405 8606 444807 8608
rect 324405 8603 324471 8606
rect 444741 8603 444807 8606
rect 56041 8530 56107 8533
rect 95141 8530 95207 8533
rect 56041 8528 95207 8530
rect 56041 8472 56046 8528
rect 56102 8472 95146 8528
rect 95202 8472 95207 8528
rect 56041 8470 95207 8472
rect 56041 8467 56107 8470
rect 95141 8467 95207 8470
rect 183737 8530 183803 8533
rect 313273 8530 313339 8533
rect 183737 8528 313339 8530
rect 183737 8472 183742 8528
rect 183798 8472 313278 8528
rect 313334 8472 313339 8528
rect 183737 8470 313339 8472
rect 183737 8467 183803 8470
rect 313273 8467 313339 8470
rect 59629 8394 59695 8397
rect 100753 8394 100819 8397
rect 59629 8392 100819 8394
rect 59629 8336 59634 8392
rect 59690 8336 100758 8392
rect 100814 8336 100819 8392
rect 59629 8334 100819 8336
rect 59629 8331 59695 8334
rect 100753 8331 100819 8334
rect 155401 8394 155467 8397
rect 317321 8394 317387 8397
rect 155401 8392 317387 8394
rect 155401 8336 155406 8392
rect 155462 8336 317326 8392
rect 317382 8336 317387 8392
rect 155401 8334 317387 8336
rect 155401 8331 155467 8334
rect 317321 8331 317387 8334
rect 335310 8334 336474 8394
rect 108113 8258 108179 8261
rect 131849 8258 131915 8261
rect 108113 8256 131915 8258
rect 108113 8200 108118 8256
rect 108174 8200 131854 8256
rect 131910 8200 131915 8256
rect 108113 8198 131915 8200
rect 108113 8195 108179 8198
rect 131849 8195 131915 8198
rect 104525 8122 104591 8125
rect 130285 8122 130351 8125
rect 104525 8120 130351 8122
rect 104525 8064 104530 8120
rect 104586 8064 130290 8120
rect 130346 8064 130351 8120
rect 104525 8062 130351 8064
rect 104525 8059 104591 8062
rect 130285 8059 130351 8062
rect 249977 8122 250043 8125
rect 335310 8122 335370 8334
rect 335537 8258 335603 8261
rect 336089 8260 336155 8261
rect 335854 8258 335860 8260
rect 335537 8256 335860 8258
rect 335537 8200 335542 8256
rect 335598 8200 335860 8256
rect 335537 8198 335860 8200
rect 335537 8195 335603 8198
rect 335854 8196 335860 8198
rect 335924 8196 335930 8260
rect 336038 8196 336044 8260
rect 336108 8258 336155 8260
rect 336414 8258 336474 8334
rect 338113 8258 338179 8261
rect 336108 8256 336200 8258
rect 336150 8200 336200 8256
rect 336108 8198 336200 8200
rect 336414 8256 338179 8258
rect 336414 8200 338118 8256
rect 338174 8200 338179 8256
rect 336414 8198 338179 8200
rect 336108 8196 336155 8198
rect 336089 8195 336155 8196
rect 338113 8195 338179 8198
rect 249977 8120 335370 8122
rect 249977 8064 249982 8120
rect 250038 8064 335370 8120
rect 249977 8062 335370 8064
rect 335721 8122 335787 8125
rect 336222 8122 336228 8124
rect 335721 8120 336228 8122
rect 335721 8064 335726 8120
rect 335782 8064 336228 8120
rect 335721 8062 336228 8064
rect 249977 8059 250043 8062
rect 335721 8059 335787 8062
rect 336222 8060 336228 8062
rect 336292 8060 336298 8124
rect 54937 7986 55003 7989
rect 86861 7986 86927 7989
rect 54937 7984 86927 7986
rect 54937 7928 54942 7984
rect 54998 7928 86866 7984
rect 86922 7928 86927 7984
rect 54937 7926 86927 7928
rect 54937 7923 55003 7926
rect 86861 7923 86927 7926
rect 87045 7986 87111 7989
rect 122465 7986 122531 7989
rect 87045 7984 122531 7986
rect 87045 7928 87050 7984
rect 87106 7928 122470 7984
rect 122526 7928 122531 7984
rect 87045 7926 122531 7928
rect 87045 7923 87111 7926
rect 122465 7923 122531 7926
rect 242893 7986 242959 7989
rect 337009 7986 337075 7989
rect 242893 7984 337075 7986
rect 242893 7928 242898 7984
rect 242954 7928 337014 7984
rect 337070 7928 337075 7984
rect 242893 7926 337075 7928
rect 242893 7923 242959 7926
rect 337009 7923 337075 7926
rect 77334 7788 77340 7852
rect 77404 7850 77410 7852
rect 83089 7850 83155 7853
rect 77404 7848 83155 7850
rect 77404 7792 83094 7848
rect 83150 7792 83155 7848
rect 77404 7790 83155 7792
rect 77404 7788 77410 7790
rect 83089 7787 83155 7790
rect 83273 7850 83339 7853
rect 120901 7850 120967 7853
rect 83273 7848 120967 7850
rect 83273 7792 83278 7848
rect 83334 7792 120906 7848
rect 120962 7792 120967 7848
rect 83273 7790 120967 7792
rect 83273 7787 83339 7790
rect 120901 7787 120967 7790
rect 239305 7850 239371 7853
rect 337285 7850 337351 7853
rect 239305 7848 337351 7850
rect 239305 7792 239310 7848
rect 239366 7792 337290 7848
rect 337346 7792 337351 7848
rect 239305 7790 337351 7792
rect 239305 7787 239371 7790
rect 337285 7787 337351 7790
rect 79685 7714 79751 7717
rect 119337 7714 119403 7717
rect 79685 7712 119403 7714
rect 79685 7656 79690 7712
rect 79746 7656 119342 7712
rect 119398 7656 119403 7712
rect 79685 7654 119403 7656
rect 79685 7651 79751 7654
rect 119337 7651 119403 7654
rect 154205 7714 154271 7717
rect 189717 7714 189783 7717
rect 154205 7712 189783 7714
rect 154205 7656 154210 7712
rect 154266 7656 189722 7712
rect 189778 7656 189783 7712
rect 154205 7654 189783 7656
rect 154205 7651 154271 7654
rect 189717 7651 189783 7654
rect 235809 7714 235875 7717
rect 337469 7714 337535 7717
rect 235809 7712 337535 7714
rect 235809 7656 235814 7712
rect 235870 7656 337474 7712
rect 337530 7656 337535 7712
rect 235809 7654 337535 7656
rect 235809 7651 235875 7654
rect 337469 7651 337535 7654
rect 72601 7578 72667 7581
rect 116209 7578 116275 7581
rect 72601 7576 116275 7578
rect 72601 7520 72606 7576
rect 72662 7520 116214 7576
rect 116270 7520 116275 7576
rect 72601 7518 116275 7520
rect 72601 7515 72667 7518
rect 116209 7515 116275 7518
rect 169569 7578 169635 7581
rect 336273 7578 336339 7581
rect 169569 7576 336339 7578
rect 169569 7520 169574 7576
rect 169630 7520 336278 7576
rect 336334 7520 336339 7576
rect 169569 7518 336339 7520
rect 169569 7515 169635 7518
rect 336273 7515 336339 7518
rect 51349 7442 51415 7445
rect 82813 7442 82879 7445
rect 51349 7440 82879 7442
rect 51349 7384 51354 7440
rect 51410 7384 82818 7440
rect 82874 7384 82879 7440
rect 51349 7382 82879 7384
rect 51349 7379 51415 7382
rect 82813 7379 82879 7382
rect 83089 7442 83155 7445
rect 98545 7442 98611 7445
rect 83089 7440 98611 7442
rect 83089 7384 83094 7440
rect 83150 7384 98550 7440
rect 98606 7384 98611 7440
rect 83089 7382 98611 7384
rect 83089 7379 83155 7382
rect 98545 7379 98611 7382
rect 98678 7380 98684 7444
rect 98748 7442 98754 7444
rect 104801 7442 104867 7445
rect 98748 7440 104867 7442
rect 98748 7384 104806 7440
rect 104862 7384 104867 7440
rect 98748 7382 104867 7384
rect 98748 7380 98754 7382
rect 104801 7379 104867 7382
rect 111609 7442 111675 7445
rect 133413 7442 133479 7445
rect 111609 7440 133479 7442
rect 111609 7384 111614 7440
rect 111670 7384 133418 7440
rect 133474 7384 133479 7440
rect 111609 7382 133479 7384
rect 111609 7379 111675 7382
rect 133413 7379 133479 7382
rect 180241 7442 180307 7445
rect 181069 7442 181135 7445
rect 193070 7442 193076 7444
rect 180241 7440 180994 7442
rect 180241 7384 180246 7440
rect 180302 7384 180994 7440
rect 180241 7382 180994 7384
rect 180241 7379 180307 7382
rect 65517 7306 65583 7309
rect 110413 7306 110479 7309
rect 65517 7304 110479 7306
rect 65517 7248 65522 7304
rect 65578 7248 110418 7304
rect 110474 7248 110479 7304
rect 65517 7246 110479 7248
rect 65517 7243 65583 7246
rect 110413 7243 110479 7246
rect 173750 7244 173756 7308
rect 173820 7306 173826 7308
rect 180793 7306 180859 7309
rect 173820 7304 180859 7306
rect 173820 7248 180798 7304
rect 180854 7248 180859 7304
rect 173820 7246 180859 7248
rect 180934 7306 180994 7382
rect 181069 7440 193076 7442
rect 181069 7384 181074 7440
rect 181130 7384 193076 7440
rect 181069 7382 193076 7384
rect 181069 7379 181135 7382
rect 193070 7380 193076 7382
rect 193140 7380 193146 7444
rect 202822 7380 202828 7444
rect 202892 7442 202898 7444
rect 212758 7442 212764 7444
rect 202892 7382 212764 7442
rect 202892 7380 202898 7382
rect 212758 7380 212764 7382
rect 212828 7380 212834 7444
rect 222837 7442 222903 7445
rect 243353 7442 243419 7445
rect 219390 7382 222762 7442
rect 219390 7306 219450 7382
rect 222702 7306 222762 7382
rect 222837 7440 243419 7442
rect 222837 7384 222842 7440
rect 222898 7384 243358 7440
rect 243414 7384 243419 7440
rect 222837 7382 243419 7384
rect 222837 7379 222903 7382
rect 243353 7379 243419 7382
rect 243486 7380 243492 7444
rect 243556 7442 243562 7444
rect 251081 7442 251147 7445
rect 256693 7442 256759 7445
rect 243556 7440 251147 7442
rect 243556 7384 251086 7440
rect 251142 7384 251147 7440
rect 243556 7382 251147 7384
rect 243556 7380 243562 7382
rect 251081 7379 251147 7382
rect 253246 7440 256759 7442
rect 253246 7384 256698 7440
rect 256754 7384 256759 7440
rect 253246 7382 256759 7384
rect 253246 7306 253306 7382
rect 256693 7379 256759 7382
rect 257061 7442 257127 7445
rect 336181 7442 336247 7445
rect 257061 7440 336247 7442
rect 257061 7384 257066 7440
rect 257122 7384 336186 7440
rect 336242 7384 336247 7440
rect 257061 7382 336247 7384
rect 257061 7379 257127 7382
rect 336181 7379 336247 7382
rect 180934 7246 219450 7306
rect 221782 7246 222578 7306
rect 222702 7246 253306 7306
rect 253473 7306 253539 7309
rect 263777 7306 263843 7309
rect 253473 7304 263843 7306
rect 253473 7248 253478 7304
rect 253534 7248 263782 7304
rect 263838 7248 263843 7304
rect 253473 7246 263843 7248
rect 173820 7244 173826 7246
rect 180793 7243 180859 7246
rect 58433 7170 58499 7173
rect 98678 7170 98684 7172
rect 58433 7168 98684 7170
rect 58433 7112 58438 7168
rect 58494 7112 98684 7168
rect 58433 7110 98684 7112
rect 58433 7107 58499 7110
rect 98678 7108 98684 7110
rect 98748 7108 98754 7172
rect 98821 7170 98887 7173
rect 114870 7170 114876 7172
rect 98821 7168 114876 7170
rect 98821 7112 98826 7168
rect 98882 7112 114876 7168
rect 98821 7110 114876 7112
rect 98821 7107 98887 7110
rect 114870 7108 114876 7110
rect 114940 7108 114946 7172
rect 166073 7170 166139 7173
rect 221782 7170 221842 7246
rect 222518 7170 222578 7246
rect 253473 7243 253539 7246
rect 263777 7243 263843 7246
rect 265617 7306 265683 7309
rect 275277 7306 275343 7309
rect 265617 7304 275343 7306
rect 265617 7248 265622 7304
rect 265678 7248 275282 7304
rect 275338 7248 275343 7304
rect 265617 7246 275343 7248
rect 265617 7243 265683 7246
rect 275277 7243 275343 7246
rect 284937 7306 285003 7309
rect 294597 7306 294663 7309
rect 284937 7304 294663 7306
rect 284937 7248 284942 7304
rect 284998 7248 294602 7304
rect 294658 7248 294663 7304
rect 284937 7246 294663 7248
rect 284937 7243 285003 7246
rect 294597 7243 294663 7246
rect 323577 7306 323643 7309
rect 336406 7306 336412 7308
rect 323577 7304 336412 7306
rect 323577 7248 323582 7304
rect 323638 7248 336412 7304
rect 323577 7246 336412 7248
rect 323577 7243 323643 7246
rect 336406 7244 336412 7246
rect 336476 7244 336482 7308
rect 243486 7170 243492 7172
rect 166073 7168 221842 7170
rect 166073 7112 166078 7168
rect 166134 7112 221842 7168
rect 166073 7110 221842 7112
rect 221966 7110 222394 7170
rect 222518 7110 243492 7170
rect 166073 7107 166139 7110
rect 62021 7034 62087 7037
rect 107653 7034 107719 7037
rect 62021 7032 107719 7034
rect 62021 6976 62026 7032
rect 62082 6976 107658 7032
rect 107714 6976 107719 7032
rect 62021 6974 107719 6976
rect 62021 6971 62087 6974
rect 107653 6971 107719 6974
rect 162485 7034 162551 7037
rect 221966 7034 222026 7110
rect 162485 7032 222026 7034
rect 162485 6976 162490 7032
rect 162546 6976 222026 7032
rect 162485 6974 222026 6976
rect 222101 7034 222167 7037
rect 222334 7034 222394 7110
rect 243486 7108 243492 7110
rect 243556 7108 243562 7172
rect 243629 7170 243695 7173
rect 264053 7170 264119 7173
rect 273161 7170 273227 7173
rect 243629 7168 258090 7170
rect 243629 7112 243634 7168
rect 243690 7112 258090 7168
rect 243629 7110 258090 7112
rect 243629 7107 243695 7110
rect 253197 7034 253263 7037
rect 222101 7032 222210 7034
rect 222101 6976 222106 7032
rect 222162 6976 222210 7032
rect 162485 6971 162551 6974
rect 222101 6971 222210 6976
rect 222334 7032 253263 7034
rect 222334 6976 253202 7032
rect 253258 6976 253263 7032
rect 222334 6974 253263 6976
rect 258030 7034 258090 7110
rect 264053 7168 273227 7170
rect 264053 7112 264058 7168
rect 264114 7112 273166 7168
rect 273222 7112 273227 7168
rect 264053 7110 273227 7112
rect 264053 7107 264119 7110
rect 273161 7107 273227 7110
rect 273437 7170 273503 7173
rect 282913 7170 282979 7173
rect 273437 7168 282979 7170
rect 273437 7112 273442 7168
rect 273498 7112 282918 7168
rect 282974 7112 282979 7168
rect 273437 7110 282979 7112
rect 273437 7107 273503 7110
rect 282913 7107 282979 7110
rect 283189 7170 283255 7173
rect 292665 7170 292731 7173
rect 283189 7168 292731 7170
rect 283189 7112 283194 7168
rect 283250 7112 292670 7168
rect 292726 7112 292731 7168
rect 283189 7110 292731 7112
rect 283189 7107 283255 7110
rect 292665 7107 292731 7110
rect 292941 7170 293007 7173
rect 321553 7170 321619 7173
rect 292941 7168 321619 7170
rect 292941 7112 292946 7168
rect 293002 7112 321558 7168
rect 321614 7112 321619 7168
rect 292941 7110 321619 7112
rect 292941 7107 293007 7110
rect 321553 7107 321619 7110
rect 321829 7170 321895 7173
rect 336365 7170 336431 7173
rect 321829 7168 336431 7170
rect 321829 7112 321834 7168
rect 321890 7112 336370 7168
rect 336426 7112 336431 7168
rect 321829 7110 336431 7112
rect 321829 7107 321895 7110
rect 336365 7107 336431 7110
rect 265617 7034 265683 7037
rect 258030 7032 265683 7034
rect 258030 6976 265622 7032
rect 265678 6976 265683 7032
rect 258030 6974 265683 6976
rect 253197 6971 253263 6974
rect 265617 6971 265683 6974
rect 275277 7034 275343 7037
rect 284937 7034 285003 7037
rect 275277 7032 285003 7034
rect 275277 6976 275282 7032
rect 275338 6976 284942 7032
rect 284998 6976 285003 7032
rect 275277 6974 285003 6976
rect 275277 6971 275343 6974
rect 284937 6971 285003 6974
rect 294597 7034 294663 7037
rect 323577 7034 323643 7037
rect 294597 7032 323643 7034
rect 294597 6976 294602 7032
rect 294658 6976 323582 7032
rect 323638 6976 323643 7032
rect 294597 6974 323643 6976
rect 294597 6971 294663 6974
rect 323577 6971 323643 6974
rect 47853 6898 47919 6901
rect 105261 6898 105327 6901
rect 47853 6896 105327 6898
rect 47853 6840 47858 6896
rect 47914 6840 105266 6896
rect 105322 6840 105327 6896
rect 47853 6838 105327 6840
rect 47853 6835 47919 6838
rect 105261 6835 105327 6838
rect 106917 6898 106983 6901
rect 192201 6898 192267 6901
rect 106917 6896 192267 6898
rect 106917 6840 106922 6896
rect 106978 6840 192206 6896
rect 192262 6840 192267 6896
rect 106917 6838 192267 6840
rect 106917 6835 106983 6838
rect 192201 6835 192267 6838
rect 193070 6836 193076 6900
rect 193140 6898 193146 6900
rect 202638 6898 202644 6900
rect 193140 6838 202644 6898
rect 193140 6836 193146 6838
rect 202638 6836 202644 6838
rect 202708 6836 202714 6900
rect 212758 6836 212764 6900
rect 212828 6898 212834 6900
rect 222150 6898 222210 6971
rect 212828 6838 222210 6898
rect 228725 6898 228791 6901
rect 337101 6898 337167 6901
rect 228725 6896 337167 6898
rect 228725 6840 228730 6896
rect 228786 6840 337106 6896
rect 337162 6840 337167 6896
rect 228725 6838 337167 6840
rect 212828 6836 212834 6838
rect 228725 6835 228791 6838
rect 337101 6835 337167 6838
rect 7649 6762 7715 6765
rect 89621 6762 89687 6765
rect 7649 6760 89687 6762
rect 7649 6704 7654 6760
rect 7710 6704 89626 6760
rect 89682 6704 89687 6760
rect 7649 6702 89687 6704
rect 7649 6699 7715 6702
rect 89621 6699 89687 6702
rect 92749 6762 92815 6765
rect 221549 6762 221615 6765
rect 336774 6762 336780 6764
rect 92749 6760 190470 6762
rect 92749 6704 92754 6760
rect 92810 6704 190470 6760
rect 92749 6702 190470 6704
rect 92749 6699 92815 6702
rect 1669 6626 1735 6629
rect 83365 6626 83431 6629
rect 1669 6624 83431 6626
rect -960 6340 480 6580
rect 1669 6568 1674 6624
rect 1730 6568 83370 6624
rect 83426 6568 83431 6624
rect 1669 6566 83431 6568
rect 1669 6563 1735 6566
rect 83365 6563 83431 6566
rect 89161 6626 89227 6629
rect 190410 6626 190470 6702
rect 221549 6760 336780 6762
rect 221549 6704 221554 6760
rect 221610 6704 336780 6760
rect 221549 6702 336780 6704
rect 221549 6699 221615 6702
rect 336774 6700 336780 6702
rect 336844 6700 336850 6764
rect 192385 6626 192451 6629
rect 89161 6624 180810 6626
rect 89161 6568 89166 6624
rect 89222 6568 180810 6624
rect 89161 6566 180810 6568
rect 190410 6624 192451 6626
rect 190410 6568 192390 6624
rect 192446 6568 192451 6624
rect 190410 6566 192451 6568
rect 89161 6563 89227 6566
rect 73797 6490 73863 6493
rect 166257 6490 166323 6493
rect 73797 6488 166323 6490
rect 73797 6432 73802 6488
rect 73858 6432 166262 6488
rect 166318 6432 166323 6488
rect 73797 6430 166323 6432
rect 180750 6490 180810 6566
rect 192385 6563 192451 6566
rect 214465 6626 214531 6629
rect 337193 6626 337259 6629
rect 214465 6624 337259 6626
rect 214465 6568 214470 6624
rect 214526 6568 337198 6624
rect 337254 6568 337259 6624
rect 214465 6566 337259 6568
rect 214465 6563 214531 6566
rect 337193 6563 337259 6566
rect 185577 6490 185643 6493
rect 180750 6488 185643 6490
rect 180750 6432 185582 6488
rect 185638 6432 185643 6488
rect 180750 6430 185643 6432
rect 73797 6427 73863 6430
rect 166257 6427 166323 6430
rect 185577 6427 185643 6430
rect 186129 6490 186195 6493
rect 338481 6490 338547 6493
rect 186129 6488 338547 6490
rect 186129 6432 186134 6488
rect 186190 6432 338486 6488
rect 338542 6432 338547 6488
rect 583520 6476 584960 6716
rect 186129 6430 338547 6432
rect 186129 6427 186195 6430
rect 338481 6427 338547 6430
rect 52545 6354 52611 6357
rect 156873 6354 156939 6357
rect 52545 6352 156939 6354
rect 52545 6296 52550 6352
rect 52606 6296 156878 6352
rect 156934 6296 156939 6352
rect 52545 6294 156939 6296
rect 52545 6291 52611 6294
rect 156873 6291 156939 6294
rect 160093 6354 160159 6357
rect 179229 6354 179295 6357
rect 160093 6352 179295 6354
rect 160093 6296 160098 6352
rect 160154 6296 179234 6352
rect 179290 6296 179295 6352
rect 160093 6294 179295 6296
rect 160093 6291 160159 6294
rect 179229 6291 179295 6294
rect 182541 6354 182607 6357
rect 338757 6354 338823 6357
rect 182541 6352 338823 6354
rect 182541 6296 182546 6352
rect 182602 6296 338762 6352
rect 338818 6296 338823 6352
rect 182541 6294 338823 6296
rect 182541 6291 182607 6294
rect 338757 6291 338823 6294
rect 13537 6218 13603 6221
rect 141233 6218 141299 6221
rect 13537 6216 141299 6218
rect 13537 6160 13542 6216
rect 13598 6160 141238 6216
rect 141294 6160 141299 6216
rect 13537 6158 141299 6160
rect 13537 6155 13603 6158
rect 141233 6155 141299 6158
rect 175457 6218 175523 6221
rect 338205 6218 338271 6221
rect 175457 6216 338271 6218
rect 175457 6160 175462 6216
rect 175518 6160 338210 6216
rect 338266 6160 338271 6216
rect 175457 6158 338271 6160
rect 175457 6155 175523 6158
rect 338205 6155 338271 6158
rect 77150 6020 77156 6084
rect 77220 6020 77226 6084
rect 117773 6082 117839 6085
rect 84150 6080 117839 6082
rect 84150 6024 117778 6080
rect 117834 6024 117839 6080
rect 84150 6022 117839 6024
rect 70342 5884 70348 5948
rect 70412 5946 70418 5948
rect 77158 5946 77218 6020
rect 70412 5886 77218 5946
rect 70412 5884 70418 5886
rect 9949 5810 10015 5813
rect 77201 5810 77267 5813
rect 9949 5808 77267 5810
rect 9949 5752 9954 5808
rect 10010 5752 77206 5808
rect 77262 5752 77267 5808
rect 9949 5750 77267 5752
rect 9949 5747 10015 5750
rect 77201 5747 77267 5750
rect 565 5674 631 5677
rect 73153 5674 73219 5677
rect 565 5672 73219 5674
rect 565 5616 570 5672
rect 626 5616 73158 5672
rect 73214 5616 73219 5672
rect 565 5614 73219 5616
rect 565 5611 631 5614
rect 73153 5611 73219 5614
rect 76189 5674 76255 5677
rect 84150 5674 84210 6022
rect 117773 6019 117839 6022
rect 185577 6082 185643 6085
rect 192477 6082 192543 6085
rect 185577 6080 192543 6082
rect 185577 6024 185582 6080
rect 185638 6024 192482 6080
rect 192538 6024 192543 6080
rect 185577 6022 192543 6024
rect 185577 6019 185643 6022
rect 192477 6019 192543 6022
rect 232221 6082 232287 6085
rect 336917 6082 336983 6085
rect 232221 6080 336983 6082
rect 232221 6024 232226 6080
rect 232282 6024 336922 6080
rect 336978 6024 336983 6080
rect 232221 6022 336983 6024
rect 232221 6019 232287 6022
rect 336917 6019 336983 6022
rect 179045 5810 179111 5813
rect 191782 5810 191788 5812
rect 179045 5808 191788 5810
rect 179045 5752 179050 5808
rect 179106 5752 191788 5808
rect 179045 5750 191788 5752
rect 179045 5747 179111 5750
rect 191782 5748 191788 5750
rect 191852 5748 191858 5812
rect 76189 5672 84210 5674
rect 76189 5616 76194 5672
rect 76250 5616 84210 5672
rect 76189 5614 84210 5616
rect 157793 5674 157859 5677
rect 185669 5674 185735 5677
rect 157793 5672 185735 5674
rect 157793 5616 157798 5672
rect 157854 5616 185674 5672
rect 185730 5616 185735 5672
rect 157793 5614 185735 5616
rect 76189 5611 76255 5614
rect 157793 5611 157859 5614
rect 185669 5611 185735 5614
rect 37181 5538 37247 5541
rect 100569 5538 100635 5541
rect 37181 5536 100635 5538
rect 37181 5480 37186 5536
rect 37242 5480 100574 5536
rect 100630 5480 100635 5536
rect 37181 5478 100635 5480
rect 37181 5475 37247 5478
rect 100569 5475 100635 5478
rect 122281 5538 122347 5541
rect 138105 5538 138171 5541
rect 122281 5536 138171 5538
rect 122281 5480 122286 5536
rect 122342 5480 138110 5536
rect 138166 5480 138171 5536
rect 122281 5478 138171 5480
rect 122281 5475 122347 5478
rect 138105 5475 138171 5478
rect 167177 5538 167243 5541
rect 180057 5538 180123 5541
rect 192109 5540 192175 5541
rect 192109 5538 192156 5540
rect 167177 5536 180123 5538
rect 167177 5480 167182 5536
rect 167238 5480 180062 5536
rect 180118 5480 180123 5536
rect 167177 5478 180123 5480
rect 192064 5536 192156 5538
rect 192064 5480 192114 5536
rect 192064 5478 192156 5480
rect 167177 5475 167243 5478
rect 180057 5475 180123 5478
rect 192109 5476 192156 5478
rect 192220 5476 192226 5540
rect 200297 5538 200363 5541
rect 338849 5538 338915 5541
rect 200297 5536 338915 5538
rect 200297 5480 200302 5536
rect 200358 5480 338854 5536
rect 338910 5480 338915 5536
rect 200297 5478 338915 5480
rect 192109 5475 192175 5476
rect 200297 5475 200363 5478
rect 338849 5475 338915 5478
rect 33593 5402 33659 5405
rect 99005 5402 99071 5405
rect 33593 5400 99071 5402
rect 33593 5344 33598 5400
rect 33654 5344 99010 5400
rect 99066 5344 99071 5400
rect 33593 5342 99071 5344
rect 33593 5339 33659 5342
rect 99005 5339 99071 5342
rect 118785 5402 118851 5405
rect 136541 5402 136607 5405
rect 118785 5400 136607 5402
rect 118785 5344 118790 5400
rect 118846 5344 136546 5400
rect 136602 5344 136607 5400
rect 118785 5342 136607 5344
rect 118785 5339 118851 5342
rect 136541 5339 136607 5342
rect 156597 5402 156663 5405
rect 174537 5402 174603 5405
rect 156597 5400 174603 5402
rect 156597 5344 156602 5400
rect 156658 5344 174542 5400
rect 174598 5344 174603 5400
rect 156597 5342 174603 5344
rect 156597 5339 156663 5342
rect 174537 5339 174603 5342
rect 288985 5402 289051 5405
rect 429101 5402 429167 5405
rect 288985 5400 429167 5402
rect 288985 5344 288990 5400
rect 289046 5344 429106 5400
rect 429162 5344 429167 5400
rect 288985 5342 429167 5344
rect 288985 5339 289051 5342
rect 429101 5339 429167 5342
rect 30097 5266 30163 5269
rect 97441 5266 97507 5269
rect 30097 5264 97507 5266
rect 30097 5208 30102 5264
rect 30158 5208 97446 5264
rect 97502 5208 97507 5264
rect 30097 5206 97507 5208
rect 30097 5203 30163 5206
rect 97441 5203 97507 5206
rect 124673 5266 124739 5269
rect 191833 5266 191899 5269
rect 124673 5264 191899 5266
rect 124673 5208 124678 5264
rect 124734 5208 191838 5264
rect 191894 5208 191899 5264
rect 124673 5206 191899 5208
rect 124673 5203 124739 5206
rect 191833 5203 191899 5206
rect 196801 5266 196867 5269
rect 338665 5266 338731 5269
rect 196801 5264 338731 5266
rect 196801 5208 196806 5264
rect 196862 5208 338670 5264
rect 338726 5208 338731 5264
rect 196801 5206 338731 5208
rect 196801 5203 196867 5206
rect 338665 5203 338731 5206
rect 26509 5130 26575 5133
rect 95877 5130 95943 5133
rect 26509 5128 95943 5130
rect 26509 5072 26514 5128
rect 26570 5072 95882 5128
rect 95938 5072 95943 5128
rect 26509 5070 95943 5072
rect 26509 5067 26575 5070
rect 95877 5067 95943 5070
rect 121085 5130 121151 5133
rect 191925 5130 191991 5133
rect 121085 5128 191991 5130
rect 121085 5072 121090 5128
rect 121146 5072 191930 5128
rect 191986 5072 191991 5128
rect 121085 5070 191991 5072
rect 121085 5067 121151 5070
rect 191925 5067 191991 5070
rect 285397 5130 285463 5133
rect 427537 5130 427603 5133
rect 285397 5128 427603 5130
rect 285397 5072 285402 5128
rect 285458 5072 427542 5128
rect 427598 5072 427603 5128
rect 285397 5070 427603 5072
rect 285397 5067 285463 5070
rect 427537 5067 427603 5070
rect 21817 4994 21883 4997
rect 94313 4994 94379 4997
rect 21817 4992 94379 4994
rect 21817 4936 21822 4992
rect 21878 4936 94318 4992
rect 94374 4936 94379 4992
rect 21817 4934 94379 4936
rect 21817 4931 21883 4934
rect 94313 4931 94379 4934
rect 117589 4994 117655 4997
rect 192017 4994 192083 4997
rect 117589 4992 192083 4994
rect 117589 4936 117594 4992
rect 117650 4936 192022 4992
rect 192078 4936 192083 4992
rect 117589 4934 192083 4936
rect 117589 4931 117655 4934
rect 192017 4931 192083 4934
rect 281901 4994 281967 4997
rect 425973 4994 426039 4997
rect 281901 4992 426039 4994
rect 281901 4936 281906 4992
rect 281962 4936 425978 4992
rect 426034 4936 426039 4992
rect 281901 4934 426039 4936
rect 281901 4931 281967 4934
rect 425973 4931 426039 4934
rect 17033 4858 17099 4861
rect 92657 4858 92723 4861
rect 17033 4856 92723 4858
rect 17033 4800 17038 4856
rect 17094 4800 92662 4856
rect 92718 4800 92723 4856
rect 17033 4798 92723 4800
rect 17033 4795 17099 4798
rect 92657 4795 92723 4798
rect 115197 4858 115263 4861
rect 134977 4858 135043 4861
rect 115197 4856 135043 4858
rect 115197 4800 115202 4856
rect 115258 4800 134982 4856
rect 135038 4800 135043 4856
rect 115197 4798 135043 4800
rect 115197 4795 115263 4798
rect 134977 4795 135043 4798
rect 163681 4858 163747 4861
rect 311433 4858 311499 4861
rect 163681 4856 311499 4858
rect 163681 4800 163686 4856
rect 163742 4800 311438 4856
rect 311494 4800 311499 4856
rect 163681 4798 311499 4800
rect 163681 4795 163747 4798
rect 311433 4795 311499 4798
rect 331581 4858 331647 4861
rect 447869 4858 447935 4861
rect 331581 4856 447935 4858
rect 331581 4800 331586 4856
rect 331642 4800 447874 4856
rect 447930 4800 447935 4856
rect 331581 4798 447935 4800
rect 331581 4795 331647 4798
rect 447869 4795 447935 4798
rect 40769 4722 40835 4725
rect 102133 4722 102199 4725
rect 40769 4720 102199 4722
rect 40769 4664 40774 4720
rect 40830 4664 102138 4720
rect 102194 4664 102199 4720
rect 40769 4662 102199 4664
rect 40769 4659 40835 4662
rect 102133 4659 102199 4662
rect 170765 4722 170831 4725
rect 178953 4722 179019 4725
rect 170765 4720 179019 4722
rect 170765 4664 170770 4720
rect 170826 4664 178958 4720
rect 179014 4664 179019 4720
rect 170765 4662 179019 4664
rect 170765 4659 170831 4662
rect 178953 4659 179019 4662
rect 306741 4722 306807 4725
rect 436921 4722 436987 4725
rect 306741 4720 436987 4722
rect 306741 4664 306746 4720
rect 306802 4664 436926 4720
rect 436982 4664 436987 4720
rect 306741 4662 436987 4664
rect 306741 4659 306807 4662
rect 436921 4659 436987 4662
rect 176653 4450 176719 4453
rect 208577 4450 208643 4453
rect 288433 4450 288499 4453
rect 176653 4448 190470 4450
rect 176653 4392 176658 4448
rect 176714 4392 190470 4448
rect 176653 4390 190470 4392
rect 176653 4387 176719 4390
rect 172973 4314 173039 4317
rect 172973 4312 177498 4314
rect 172973 4256 172978 4312
rect 173034 4256 177498 4312
rect 172973 4254 177498 4256
rect 172973 4251 173039 4254
rect 8753 4178 8819 4181
rect 40677 4178 40743 4181
rect 8753 4176 40743 4178
rect 8753 4120 8758 4176
rect 8814 4120 40682 4176
rect 40738 4120 40743 4176
rect 8753 4118 40743 4120
rect 8753 4115 8819 4118
rect 40677 4115 40743 4118
rect 174261 4178 174327 4181
rect 177246 4178 177252 4180
rect 174261 4176 177252 4178
rect 174261 4120 174266 4176
rect 174322 4120 177252 4176
rect 174261 4118 177252 4120
rect 174261 4115 174327 4118
rect 177246 4116 177252 4118
rect 177316 4116 177322 4180
rect 177438 4178 177498 4254
rect 189390 4178 189396 4180
rect 177438 4118 189396 4178
rect 189390 4116 189396 4118
rect 189460 4116 189466 4180
rect 190410 4178 190470 4390
rect 208577 4448 288499 4450
rect 208577 4392 208582 4448
rect 208638 4392 288438 4448
rect 288494 4392 288499 4448
rect 208577 4390 288499 4392
rect 208577 4387 208643 4390
rect 288433 4387 288499 4390
rect 201493 4314 201559 4317
rect 285581 4314 285647 4317
rect 201493 4312 285647 4314
rect 201493 4256 201498 4312
rect 201554 4256 285586 4312
rect 285642 4256 285647 4312
rect 201493 4254 285647 4256
rect 201493 4251 201559 4254
rect 285581 4251 285647 4254
rect 307661 4178 307727 4181
rect 190410 4176 307727 4178
rect 190410 4120 307666 4176
rect 307722 4120 307727 4176
rect 190410 4118 307727 4120
rect 307661 4115 307727 4118
rect 335169 4178 335235 4181
rect 344921 4178 344987 4181
rect 335169 4176 344987 4178
rect 335169 4120 335174 4176
rect 335230 4120 344926 4176
rect 344982 4120 344987 4176
rect 335169 4118 344987 4120
rect 335169 4115 335235 4118
rect 344921 4115 344987 4118
rect 40677 4042 40743 4045
rect 26190 4040 40743 4042
rect 26190 3984 40682 4040
rect 40738 3984 40743 4040
rect 26190 3982 40743 3984
rect 6453 3770 6519 3773
rect 26190 3770 26250 3982
rect 40677 3979 40743 3982
rect 99833 4042 99899 4045
rect 190453 4042 190519 4045
rect 99833 4040 190519 4042
rect 99833 3984 99838 4040
rect 99894 3984 190458 4040
rect 190514 3984 190519 4040
rect 99833 3982 190519 3984
rect 99833 3979 99899 3982
rect 190453 3979 190519 3982
rect 190821 4042 190887 4045
rect 191046 4042 191052 4044
rect 190821 4040 191052 4042
rect 190821 3984 190826 4040
rect 190882 3984 191052 4040
rect 190821 3982 191052 3984
rect 190821 3979 190887 3982
rect 191046 3980 191052 3982
rect 191116 3980 191122 4044
rect 193213 4042 193279 4045
rect 338481 4042 338547 4045
rect 193213 4040 338547 4042
rect 193213 3984 193218 4040
rect 193274 3984 338486 4040
rect 338542 3984 338547 4040
rect 193213 3982 338547 3984
rect 193213 3979 193279 3982
rect 338481 3979 338547 3982
rect 338665 4042 338731 4045
rect 349705 4042 349771 4045
rect 356145 4042 356211 4045
rect 338665 4040 349771 4042
rect 338665 3984 338670 4040
rect 338726 3984 349710 4040
rect 349766 3984 349771 4040
rect 338665 3982 349771 3984
rect 338665 3979 338731 3982
rect 349705 3979 349771 3982
rect 349846 4040 356211 4042
rect 349846 3984 356150 4040
rect 356206 3984 356211 4040
rect 349846 3982 356211 3984
rect 35985 3906 36051 3909
rect 89713 3906 89779 3909
rect 172973 3906 173039 3909
rect 35985 3904 89779 3906
rect 35985 3848 35990 3904
rect 36046 3848 89718 3904
rect 89774 3848 89779 3904
rect 35985 3846 89779 3848
rect 35985 3843 36051 3846
rect 89713 3843 89779 3846
rect 93810 3904 173039 3906
rect 93810 3848 172978 3904
rect 173034 3848 173039 3904
rect 93810 3846 173039 3848
rect 93810 3770 93870 3846
rect 172973 3843 173039 3846
rect 173157 3906 173223 3909
rect 173382 3906 173388 3908
rect 173157 3904 173388 3906
rect 173157 3848 173162 3904
rect 173218 3848 173388 3904
rect 173157 3846 173388 3848
rect 173157 3843 173223 3846
rect 173382 3844 173388 3846
rect 173452 3844 173458 3908
rect 173617 3906 173683 3909
rect 173617 3904 335370 3906
rect 173617 3848 173622 3904
rect 173678 3848 335370 3904
rect 173617 3846 335370 3848
rect 173617 3843 173683 3846
rect 6453 3768 26250 3770
rect 6453 3712 6458 3768
rect 6514 3712 26250 3768
rect 6453 3710 26250 3712
rect 35850 3710 93870 3770
rect 6453 3707 6519 3710
rect 24209 3634 24275 3637
rect 35850 3634 35910 3710
rect 94998 3708 95004 3772
rect 95068 3770 95074 3772
rect 95141 3770 95207 3773
rect 95068 3768 95207 3770
rect 95068 3712 95146 3768
rect 95202 3712 95207 3768
rect 95068 3710 95207 3712
rect 95068 3708 95074 3710
rect 95141 3707 95207 3710
rect 96245 3770 96311 3773
rect 190545 3770 190611 3773
rect 96245 3768 190611 3770
rect 96245 3712 96250 3768
rect 96306 3712 190550 3768
rect 190606 3712 190611 3768
rect 96245 3710 190611 3712
rect 96245 3707 96311 3710
rect 190545 3707 190611 3710
rect 205081 3770 205147 3773
rect 233233 3770 233299 3773
rect 205081 3768 233299 3770
rect 205081 3712 205086 3768
rect 205142 3712 233238 3768
rect 233294 3712 233299 3768
rect 205081 3710 233299 3712
rect 205081 3707 205147 3710
rect 233233 3707 233299 3710
rect 233417 3770 233483 3773
rect 243537 3770 243603 3773
rect 233417 3768 243603 3770
rect 233417 3712 233422 3768
rect 233478 3712 243542 3768
rect 243598 3712 243603 3768
rect 233417 3710 243603 3712
rect 233417 3707 233483 3710
rect 243537 3707 243603 3710
rect 248321 3770 248387 3773
rect 335169 3770 335235 3773
rect 248321 3768 335235 3770
rect 248321 3712 248326 3768
rect 248382 3712 335174 3768
rect 335230 3712 335235 3768
rect 248321 3710 335235 3712
rect 335310 3770 335370 3846
rect 335486 3844 335492 3908
rect 335556 3906 335562 3908
rect 349846 3906 349906 3982
rect 356145 3979 356211 3982
rect 356329 4042 356395 4045
rect 398097 4042 398163 4045
rect 356329 4040 398163 4042
rect 356329 3984 356334 4040
rect 356390 3984 398102 4040
rect 398158 3984 398163 4040
rect 356329 3982 398163 3984
rect 356329 3979 356395 3982
rect 398097 3979 398163 3982
rect 398281 4042 398347 4045
rect 414657 4042 414723 4045
rect 398281 4040 414723 4042
rect 398281 3984 398286 4040
rect 398342 3984 414662 4040
rect 414718 3984 414723 4040
rect 398281 3982 414723 3984
rect 398281 3979 398347 3982
rect 414657 3979 414723 3982
rect 335556 3846 349906 3906
rect 349981 3906 350047 3909
rect 450997 3906 451063 3909
rect 349981 3904 451063 3906
rect 349981 3848 349986 3904
rect 350042 3848 451002 3904
rect 451058 3848 451063 3904
rect 349981 3846 451063 3848
rect 335556 3844 335562 3846
rect 349981 3843 350047 3846
rect 450997 3843 451063 3846
rect 338297 3770 338363 3773
rect 335310 3768 338363 3770
rect 335310 3712 338302 3768
rect 338358 3712 338363 3768
rect 335310 3710 338363 3712
rect 248321 3707 248387 3710
rect 335169 3707 335235 3710
rect 338297 3707 338363 3710
rect 338481 3770 338547 3773
rect 339493 3770 339559 3773
rect 338481 3768 339559 3770
rect 338481 3712 338486 3768
rect 338542 3712 339498 3768
rect 339554 3712 339559 3768
rect 338481 3710 339559 3712
rect 338481 3707 338547 3710
rect 339493 3707 339559 3710
rect 344921 3770 344987 3773
rect 409086 3770 409092 3772
rect 344921 3768 409092 3770
rect 344921 3712 344926 3768
rect 344982 3712 409092 3768
rect 344921 3710 409092 3712
rect 344921 3707 344987 3710
rect 409086 3708 409092 3710
rect 409156 3708 409162 3772
rect 24209 3632 35910 3634
rect 24209 3576 24214 3632
rect 24270 3576 35910 3632
rect 24209 3574 35910 3576
rect 40677 3634 40743 3637
rect 88057 3634 88123 3637
rect 40677 3632 88123 3634
rect 40677 3576 40682 3632
rect 40738 3576 88062 3632
rect 88118 3576 88123 3632
rect 40677 3574 88123 3576
rect 24209 3571 24275 3574
rect 40677 3571 40743 3574
rect 88057 3571 88123 3574
rect 88977 3634 89043 3637
rect 219249 3634 219315 3637
rect 411989 3634 412055 3637
rect 88977 3632 185594 3634
rect 88977 3576 88982 3632
rect 89038 3576 185594 3632
rect 88977 3574 185594 3576
rect 88977 3571 89043 3574
rect 185534 3501 185594 3574
rect 219249 3632 412055 3634
rect 219249 3576 219254 3632
rect 219310 3576 411994 3632
rect 412050 3576 412055 3632
rect 219249 3574 412055 3576
rect 219249 3571 219315 3574
rect 411989 3571 412055 3574
rect 27705 3498 27771 3501
rect 27838 3498 27844 3500
rect 27705 3496 27844 3498
rect 27705 3440 27710 3496
rect 27766 3440 27844 3496
rect 27705 3438 27844 3440
rect 27705 3435 27771 3438
rect 27838 3436 27844 3438
rect 27908 3436 27914 3500
rect 39573 3498 39639 3501
rect 39573 3496 185226 3498
rect 39573 3440 39578 3496
rect 39634 3440 185226 3496
rect 39573 3438 185226 3440
rect 185534 3496 185643 3501
rect 189533 3498 189599 3501
rect 185534 3440 185582 3496
rect 185638 3440 185643 3496
rect 185534 3438 185643 3440
rect 39573 3435 39639 3438
rect 28901 3362 28967 3365
rect 185025 3362 185091 3365
rect 28901 3360 185091 3362
rect 28901 3304 28906 3360
rect 28962 3304 185030 3360
rect 185086 3304 185091 3360
rect 28901 3302 185091 3304
rect 185166 3362 185226 3438
rect 185577 3435 185643 3438
rect 185718 3496 189599 3498
rect 185718 3440 189538 3496
rect 189594 3440 189599 3496
rect 185718 3438 189599 3440
rect 185718 3362 185778 3438
rect 189533 3435 189599 3438
rect 189717 3498 189783 3501
rect 193857 3498 193923 3501
rect 189717 3496 193923 3498
rect 189717 3440 189722 3496
rect 189778 3440 193862 3496
rect 193918 3440 193923 3496
rect 189717 3438 193923 3440
rect 189717 3435 189783 3438
rect 193857 3435 193923 3438
rect 226333 3498 226399 3501
rect 419717 3498 419783 3501
rect 226333 3496 419783 3498
rect 226333 3440 226338 3496
rect 226394 3440 419722 3496
rect 419778 3440 419783 3496
rect 226333 3438 419783 3440
rect 226333 3435 226399 3438
rect 419717 3435 419783 3438
rect 185166 3302 185778 3362
rect 212165 3362 212231 3365
rect 410374 3362 410380 3364
rect 212165 3360 410380 3362
rect 212165 3304 212170 3360
rect 212226 3304 410380 3360
rect 212165 3302 410380 3304
rect 28901 3299 28967 3302
rect 185025 3299 185091 3302
rect 212165 3299 212231 3302
rect 410374 3300 410380 3302
rect 410444 3300 410450 3364
rect 43069 3226 43135 3229
rect 44030 3226 44036 3228
rect 43069 3224 44036 3226
rect 43069 3168 43074 3224
rect 43130 3168 44036 3224
rect 43069 3166 44036 3168
rect 43069 3163 43135 3166
rect 44030 3164 44036 3166
rect 44100 3164 44106 3228
rect 57237 3226 57303 3229
rect 57830 3226 57836 3228
rect 57237 3224 57836 3226
rect 57237 3168 57242 3224
rect 57298 3168 57836 3224
rect 57237 3166 57836 3168
rect 57237 3163 57303 3166
rect 57830 3164 57836 3166
rect 57900 3164 57906 3228
rect 66713 3226 66779 3229
rect 67398 3226 67404 3228
rect 66713 3224 67404 3226
rect 66713 3168 66718 3224
rect 66774 3168 67404 3224
rect 66713 3166 67404 3168
rect 66713 3163 66779 3166
rect 67398 3164 67404 3166
rect 67468 3164 67474 3228
rect 69105 3226 69171 3229
rect 70342 3226 70348 3228
rect 69105 3224 70348 3226
rect 69105 3168 69110 3224
rect 69166 3168 70348 3224
rect 69105 3166 70348 3168
rect 69105 3163 69171 3166
rect 70342 3164 70348 3166
rect 70412 3164 70418 3228
rect 82077 3226 82143 3229
rect 88977 3226 89043 3229
rect 82077 3224 89043 3226
rect 82077 3168 82082 3224
rect 82138 3168 88982 3224
rect 89038 3168 89043 3224
rect 82077 3166 89043 3168
rect 82077 3163 82143 3166
rect 88977 3163 89043 3166
rect 103329 3226 103395 3229
rect 192293 3226 192359 3229
rect 103329 3224 192359 3226
rect 103329 3168 103334 3224
rect 103390 3168 192298 3224
rect 192354 3168 192359 3224
rect 103329 3166 192359 3168
rect 103329 3163 103395 3166
rect 192293 3163 192359 3166
rect 203885 3226 203951 3229
rect 204110 3226 204116 3228
rect 203885 3224 204116 3226
rect 203885 3168 203890 3224
rect 203946 3168 204116 3224
rect 203885 3166 204116 3168
rect 203885 3163 203951 3166
rect 204110 3164 204116 3166
rect 204180 3164 204186 3228
rect 225137 3226 225203 3229
rect 339677 3226 339743 3229
rect 225137 3224 339743 3226
rect 225137 3168 225142 3224
rect 225198 3168 339682 3224
rect 339738 3168 339743 3224
rect 225137 3166 339743 3168
rect 225137 3163 225203 3166
rect 339677 3163 339743 3166
rect 356145 3226 356211 3229
rect 398097 3226 398163 3229
rect 403617 3226 403683 3229
rect 356145 3224 393330 3226
rect 356145 3168 356150 3224
rect 356206 3168 393330 3224
rect 356145 3166 393330 3168
rect 356145 3163 356211 3166
rect 2865 3090 2931 3093
rect 81433 3090 81499 3093
rect 2865 3088 81499 3090
rect 2865 3032 2870 3088
rect 2926 3032 81438 3088
rect 81494 3032 81499 3088
rect 2865 3030 81499 3032
rect 2865 3027 2931 3030
rect 81433 3027 81499 3030
rect 171961 3090 172027 3093
rect 173617 3090 173683 3093
rect 171961 3088 173683 3090
rect 171961 3032 171966 3088
rect 172022 3032 173622 3088
rect 173678 3032 173683 3088
rect 171961 3030 173683 3032
rect 171961 3027 172027 3030
rect 173617 3027 173683 3030
rect 185577 3090 185643 3093
rect 192569 3090 192635 3093
rect 185577 3088 192635 3090
rect 185577 3032 185582 3088
rect 185638 3032 192574 3088
rect 192630 3032 192635 3088
rect 185577 3030 192635 3032
rect 185577 3027 185643 3030
rect 192569 3027 192635 3030
rect 194409 3090 194475 3093
rect 226425 3090 226491 3093
rect 194409 3088 226491 3090
rect 194409 3032 194414 3088
rect 194470 3032 226430 3088
rect 226486 3032 226491 3088
rect 194409 3030 226491 3032
rect 194409 3027 194475 3030
rect 226425 3027 226491 3030
rect 243537 3090 243603 3093
rect 335118 3090 335124 3092
rect 243537 3088 335124 3090
rect 243537 3032 243542 3088
rect 243598 3032 335124 3088
rect 243537 3030 335124 3032
rect 243537 3027 243603 3030
rect 335118 3028 335124 3030
rect 335188 3028 335194 3092
rect 393270 3090 393330 3166
rect 398097 3224 403683 3226
rect 398097 3168 398102 3224
rect 398158 3168 403622 3224
rect 403678 3168 403683 3224
rect 398097 3166 403683 3168
rect 398097 3163 398163 3166
rect 403617 3163 403683 3166
rect 398281 3090 398347 3093
rect 393270 3088 398347 3090
rect 393270 3032 398286 3088
rect 398342 3032 398347 3088
rect 393270 3030 398347 3032
rect 398281 3027 398347 3030
rect 14733 2954 14799 2957
rect 102133 2954 102199 2957
rect 14733 2952 102199 2954
rect 14733 2896 14738 2952
rect 14794 2896 102138 2952
rect 102194 2896 102199 2952
rect 14733 2894 102199 2896
rect 14733 2891 14799 2894
rect 102133 2891 102199 2894
rect 113582 2892 113588 2956
rect 113652 2954 113658 2956
rect 114001 2954 114067 2957
rect 113652 2952 114067 2954
rect 113652 2896 114006 2952
rect 114062 2896 114067 2952
rect 113652 2894 114067 2896
rect 113652 2892 113658 2894
rect 114001 2891 114067 2894
rect 185025 2954 185091 2957
rect 189625 2954 189691 2957
rect 185025 2952 189691 2954
rect 185025 2896 185030 2952
rect 185086 2896 189630 2952
rect 189686 2896 189691 2952
rect 185025 2894 189691 2896
rect 185025 2891 185091 2894
rect 189625 2891 189691 2894
rect 190821 2954 190887 2957
rect 224953 2954 225019 2957
rect 190821 2952 225019 2954
rect 190821 2896 190826 2952
rect 190882 2896 224958 2952
rect 225014 2896 225019 2952
rect 190821 2894 225019 2896
rect 190821 2891 190887 2894
rect 224953 2891 225019 2894
rect 233233 2954 233299 2957
rect 248321 2954 248387 2957
rect 233233 2952 248387 2954
rect 233233 2896 233238 2952
rect 233294 2896 248326 2952
rect 248382 2896 248387 2952
rect 233233 2894 248387 2896
rect 233233 2891 233299 2894
rect 248321 2891 248387 2894
rect 296069 2954 296135 2957
rect 296662 2954 296668 2956
rect 296069 2952 296668 2954
rect 296069 2896 296074 2952
rect 296130 2896 296668 2952
rect 296069 2894 296668 2896
rect 296069 2891 296135 2894
rect 296662 2892 296668 2894
rect 296732 2892 296738 2956
rect 12341 2820 12407 2821
rect 12341 2818 12388 2820
rect 12296 2816 12388 2818
rect 12296 2760 12346 2816
rect 12296 2758 12388 2760
rect 12341 2756 12388 2758
rect 12452 2756 12458 2820
rect 19425 2818 19491 2821
rect 172421 2818 172487 2821
rect 19425 2816 172487 2818
rect 19425 2760 19430 2816
rect 19486 2760 172426 2816
rect 172482 2760 172487 2816
rect 19425 2758 172487 2760
rect 12341 2755 12407 2756
rect 19425 2755 19491 2758
rect 172421 2755 172487 2758
rect 197905 2818 197971 2821
rect 233877 2818 233943 2821
rect 197905 2816 233943 2818
rect 197905 2760 197910 2816
rect 197966 2760 233882 2816
rect 233938 2760 233943 2816
rect 197905 2758 233943 2760
rect 197905 2755 197971 2758
rect 233877 2755 233943 2758
<< via3 >>
rect 192340 700436 192404 700500
rect 191788 177108 191852 177172
rect 191236 127060 191300 127124
rect 335860 117404 335924 117468
rect 336044 116452 336108 116516
rect 190500 114548 190564 114612
rect 338988 111692 339052 111756
rect 336780 110740 336844 110804
rect 338620 109788 338684 109852
rect 336228 107884 336292 107948
rect 338436 105980 338500 106044
rect 189396 98908 189460 98972
rect 336412 98636 336476 98700
rect 338804 98364 338868 98428
rect 190868 92652 190932 92716
rect 192340 86396 192404 86460
rect 191972 83268 192036 83332
rect 335676 81228 335740 81292
rect 335676 80548 335740 80612
rect 324268 78508 324332 78572
rect 431908 78508 431972 78572
rect 162900 78100 162964 78164
rect 145052 77828 145116 77892
rect 175228 77828 175292 77892
rect 410380 77828 410444 77892
rect 91140 77344 91204 77348
rect 91140 77288 91154 77344
rect 91154 77288 91204 77344
rect 91140 77284 91204 77288
rect 114876 77284 114940 77348
rect 409092 77284 409156 77348
rect 338620 10372 338684 10436
rect 338804 10236 338868 10300
rect 335860 8196 335924 8260
rect 336044 8256 336108 8260
rect 336044 8200 336094 8256
rect 336094 8200 336108 8256
rect 336044 8196 336108 8200
rect 336228 8060 336292 8124
rect 77340 7788 77404 7852
rect 98684 7380 98748 7444
rect 173756 7244 173820 7308
rect 193076 7380 193140 7444
rect 202828 7380 202892 7444
rect 212764 7380 212828 7444
rect 243492 7380 243556 7444
rect 98684 7108 98748 7172
rect 114876 7108 114940 7172
rect 336412 7244 336476 7308
rect 243492 7108 243556 7172
rect 193076 6836 193140 6900
rect 202644 6836 202708 6900
rect 212764 6836 212828 6900
rect 336780 6700 336844 6764
rect 77156 6020 77220 6084
rect 70348 5884 70412 5948
rect 191788 5748 191852 5812
rect 192156 5536 192220 5540
rect 192156 5480 192170 5536
rect 192170 5480 192220 5536
rect 192156 5476 192220 5480
rect 177252 4116 177316 4180
rect 189396 4116 189460 4180
rect 191052 3980 191116 4044
rect 173388 3844 173452 3908
rect 95004 3708 95068 3772
rect 335492 3844 335556 3908
rect 409092 3708 409156 3772
rect 27844 3436 27908 3500
rect 410380 3300 410444 3364
rect 44036 3164 44100 3228
rect 57836 3164 57900 3228
rect 67404 3164 67468 3228
rect 70348 3164 70412 3228
rect 204116 3164 204180 3228
rect 335124 3028 335188 3092
rect 113588 2892 113652 2956
rect 296668 2892 296732 2956
rect 12388 2816 12452 2820
rect 12388 2760 12402 2816
rect 12402 2760 12452 2816
rect 12388 2756 12452 2760
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677894 -8106 711002
rect -8726 677658 -8694 677894
rect -8458 677658 -8374 677894
rect -8138 677658 -8106 677894
rect -8726 677574 -8106 677658
rect -8726 677338 -8694 677574
rect -8458 677338 -8374 677574
rect -8138 677338 -8106 677574
rect -8726 641894 -8106 677338
rect -8726 641658 -8694 641894
rect -8458 641658 -8374 641894
rect -8138 641658 -8106 641894
rect -8726 641574 -8106 641658
rect -8726 641338 -8694 641574
rect -8458 641338 -8374 641574
rect -8138 641338 -8106 641574
rect -8726 605894 -8106 641338
rect -8726 605658 -8694 605894
rect -8458 605658 -8374 605894
rect -8138 605658 -8106 605894
rect -8726 605574 -8106 605658
rect -8726 605338 -8694 605574
rect -8458 605338 -8374 605574
rect -8138 605338 -8106 605574
rect -8726 569894 -8106 605338
rect -8726 569658 -8694 569894
rect -8458 569658 -8374 569894
rect -8138 569658 -8106 569894
rect -8726 569574 -8106 569658
rect -8726 569338 -8694 569574
rect -8458 569338 -8374 569574
rect -8138 569338 -8106 569574
rect -8726 533894 -8106 569338
rect -8726 533658 -8694 533894
rect -8458 533658 -8374 533894
rect -8138 533658 -8106 533894
rect -8726 533574 -8106 533658
rect -8726 533338 -8694 533574
rect -8458 533338 -8374 533574
rect -8138 533338 -8106 533574
rect -8726 497894 -8106 533338
rect -8726 497658 -8694 497894
rect -8458 497658 -8374 497894
rect -8138 497658 -8106 497894
rect -8726 497574 -8106 497658
rect -8726 497338 -8694 497574
rect -8458 497338 -8374 497574
rect -8138 497338 -8106 497574
rect -8726 461894 -8106 497338
rect -8726 461658 -8694 461894
rect -8458 461658 -8374 461894
rect -8138 461658 -8106 461894
rect -8726 461574 -8106 461658
rect -8726 461338 -8694 461574
rect -8458 461338 -8374 461574
rect -8138 461338 -8106 461574
rect -8726 425894 -8106 461338
rect -8726 425658 -8694 425894
rect -8458 425658 -8374 425894
rect -8138 425658 -8106 425894
rect -8726 425574 -8106 425658
rect -8726 425338 -8694 425574
rect -8458 425338 -8374 425574
rect -8138 425338 -8106 425574
rect -8726 389894 -8106 425338
rect -8726 389658 -8694 389894
rect -8458 389658 -8374 389894
rect -8138 389658 -8106 389894
rect -8726 389574 -8106 389658
rect -8726 389338 -8694 389574
rect -8458 389338 -8374 389574
rect -8138 389338 -8106 389574
rect -8726 353894 -8106 389338
rect -8726 353658 -8694 353894
rect -8458 353658 -8374 353894
rect -8138 353658 -8106 353894
rect -8726 353574 -8106 353658
rect -8726 353338 -8694 353574
rect -8458 353338 -8374 353574
rect -8138 353338 -8106 353574
rect -8726 317894 -8106 353338
rect -8726 317658 -8694 317894
rect -8458 317658 -8374 317894
rect -8138 317658 -8106 317894
rect -8726 317574 -8106 317658
rect -8726 317338 -8694 317574
rect -8458 317338 -8374 317574
rect -8138 317338 -8106 317574
rect -8726 281894 -8106 317338
rect -8726 281658 -8694 281894
rect -8458 281658 -8374 281894
rect -8138 281658 -8106 281894
rect -8726 281574 -8106 281658
rect -8726 281338 -8694 281574
rect -8458 281338 -8374 281574
rect -8138 281338 -8106 281574
rect -8726 245894 -8106 281338
rect -8726 245658 -8694 245894
rect -8458 245658 -8374 245894
rect -8138 245658 -8106 245894
rect -8726 245574 -8106 245658
rect -8726 245338 -8694 245574
rect -8458 245338 -8374 245574
rect -8138 245338 -8106 245574
rect -8726 209894 -8106 245338
rect -8726 209658 -8694 209894
rect -8458 209658 -8374 209894
rect -8138 209658 -8106 209894
rect -8726 209574 -8106 209658
rect -8726 209338 -8694 209574
rect -8458 209338 -8374 209574
rect -8138 209338 -8106 209574
rect -8726 173894 -8106 209338
rect -8726 173658 -8694 173894
rect -8458 173658 -8374 173894
rect -8138 173658 -8106 173894
rect -8726 173574 -8106 173658
rect -8726 173338 -8694 173574
rect -8458 173338 -8374 173574
rect -8138 173338 -8106 173574
rect -8726 137894 -8106 173338
rect -8726 137658 -8694 137894
rect -8458 137658 -8374 137894
rect -8138 137658 -8106 137894
rect -8726 137574 -8106 137658
rect -8726 137338 -8694 137574
rect -8458 137338 -8374 137574
rect -8138 137338 -8106 137574
rect -8726 101894 -8106 137338
rect -8726 101658 -8694 101894
rect -8458 101658 -8374 101894
rect -8138 101658 -8106 101894
rect -8726 101574 -8106 101658
rect -8726 101338 -8694 101574
rect -8458 101338 -8374 101574
rect -8138 101338 -8106 101574
rect -8726 65894 -8106 101338
rect -8726 65658 -8694 65894
rect -8458 65658 -8374 65894
rect -8138 65658 -8106 65894
rect -8726 65574 -8106 65658
rect -8726 65338 -8694 65574
rect -8458 65338 -8374 65574
rect -8138 65338 -8106 65574
rect -8726 29894 -8106 65338
rect -8726 29658 -8694 29894
rect -8458 29658 -8374 29894
rect -8138 29658 -8106 29894
rect -8726 29574 -8106 29658
rect -8726 29338 -8694 29574
rect -8458 29338 -8374 29574
rect -8138 29338 -8106 29574
rect -8726 -7066 -8106 29338
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 674174 -7146 710042
rect -7766 673938 -7734 674174
rect -7498 673938 -7414 674174
rect -7178 673938 -7146 674174
rect -7766 673854 -7146 673938
rect -7766 673618 -7734 673854
rect -7498 673618 -7414 673854
rect -7178 673618 -7146 673854
rect -7766 638174 -7146 673618
rect -7766 637938 -7734 638174
rect -7498 637938 -7414 638174
rect -7178 637938 -7146 638174
rect -7766 637854 -7146 637938
rect -7766 637618 -7734 637854
rect -7498 637618 -7414 637854
rect -7178 637618 -7146 637854
rect -7766 602174 -7146 637618
rect -7766 601938 -7734 602174
rect -7498 601938 -7414 602174
rect -7178 601938 -7146 602174
rect -7766 601854 -7146 601938
rect -7766 601618 -7734 601854
rect -7498 601618 -7414 601854
rect -7178 601618 -7146 601854
rect -7766 566174 -7146 601618
rect -7766 565938 -7734 566174
rect -7498 565938 -7414 566174
rect -7178 565938 -7146 566174
rect -7766 565854 -7146 565938
rect -7766 565618 -7734 565854
rect -7498 565618 -7414 565854
rect -7178 565618 -7146 565854
rect -7766 530174 -7146 565618
rect -7766 529938 -7734 530174
rect -7498 529938 -7414 530174
rect -7178 529938 -7146 530174
rect -7766 529854 -7146 529938
rect -7766 529618 -7734 529854
rect -7498 529618 -7414 529854
rect -7178 529618 -7146 529854
rect -7766 494174 -7146 529618
rect -7766 493938 -7734 494174
rect -7498 493938 -7414 494174
rect -7178 493938 -7146 494174
rect -7766 493854 -7146 493938
rect -7766 493618 -7734 493854
rect -7498 493618 -7414 493854
rect -7178 493618 -7146 493854
rect -7766 458174 -7146 493618
rect -7766 457938 -7734 458174
rect -7498 457938 -7414 458174
rect -7178 457938 -7146 458174
rect -7766 457854 -7146 457938
rect -7766 457618 -7734 457854
rect -7498 457618 -7414 457854
rect -7178 457618 -7146 457854
rect -7766 422174 -7146 457618
rect -7766 421938 -7734 422174
rect -7498 421938 -7414 422174
rect -7178 421938 -7146 422174
rect -7766 421854 -7146 421938
rect -7766 421618 -7734 421854
rect -7498 421618 -7414 421854
rect -7178 421618 -7146 421854
rect -7766 386174 -7146 421618
rect -7766 385938 -7734 386174
rect -7498 385938 -7414 386174
rect -7178 385938 -7146 386174
rect -7766 385854 -7146 385938
rect -7766 385618 -7734 385854
rect -7498 385618 -7414 385854
rect -7178 385618 -7146 385854
rect -7766 350174 -7146 385618
rect -7766 349938 -7734 350174
rect -7498 349938 -7414 350174
rect -7178 349938 -7146 350174
rect -7766 349854 -7146 349938
rect -7766 349618 -7734 349854
rect -7498 349618 -7414 349854
rect -7178 349618 -7146 349854
rect -7766 314174 -7146 349618
rect -7766 313938 -7734 314174
rect -7498 313938 -7414 314174
rect -7178 313938 -7146 314174
rect -7766 313854 -7146 313938
rect -7766 313618 -7734 313854
rect -7498 313618 -7414 313854
rect -7178 313618 -7146 313854
rect -7766 278174 -7146 313618
rect -7766 277938 -7734 278174
rect -7498 277938 -7414 278174
rect -7178 277938 -7146 278174
rect -7766 277854 -7146 277938
rect -7766 277618 -7734 277854
rect -7498 277618 -7414 277854
rect -7178 277618 -7146 277854
rect -7766 242174 -7146 277618
rect -7766 241938 -7734 242174
rect -7498 241938 -7414 242174
rect -7178 241938 -7146 242174
rect -7766 241854 -7146 241938
rect -7766 241618 -7734 241854
rect -7498 241618 -7414 241854
rect -7178 241618 -7146 241854
rect -7766 206174 -7146 241618
rect -7766 205938 -7734 206174
rect -7498 205938 -7414 206174
rect -7178 205938 -7146 206174
rect -7766 205854 -7146 205938
rect -7766 205618 -7734 205854
rect -7498 205618 -7414 205854
rect -7178 205618 -7146 205854
rect -7766 170174 -7146 205618
rect -7766 169938 -7734 170174
rect -7498 169938 -7414 170174
rect -7178 169938 -7146 170174
rect -7766 169854 -7146 169938
rect -7766 169618 -7734 169854
rect -7498 169618 -7414 169854
rect -7178 169618 -7146 169854
rect -7766 134174 -7146 169618
rect -7766 133938 -7734 134174
rect -7498 133938 -7414 134174
rect -7178 133938 -7146 134174
rect -7766 133854 -7146 133938
rect -7766 133618 -7734 133854
rect -7498 133618 -7414 133854
rect -7178 133618 -7146 133854
rect -7766 98174 -7146 133618
rect -7766 97938 -7734 98174
rect -7498 97938 -7414 98174
rect -7178 97938 -7146 98174
rect -7766 97854 -7146 97938
rect -7766 97618 -7734 97854
rect -7498 97618 -7414 97854
rect -7178 97618 -7146 97854
rect -7766 62174 -7146 97618
rect -7766 61938 -7734 62174
rect -7498 61938 -7414 62174
rect -7178 61938 -7146 62174
rect -7766 61854 -7146 61938
rect -7766 61618 -7734 61854
rect -7498 61618 -7414 61854
rect -7178 61618 -7146 61854
rect -7766 26174 -7146 61618
rect -7766 25938 -7734 26174
rect -7498 25938 -7414 26174
rect -7178 25938 -7146 26174
rect -7766 25854 -7146 25938
rect -7766 25618 -7734 25854
rect -7498 25618 -7414 25854
rect -7178 25618 -7146 25854
rect -7766 -6106 -7146 25618
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670454 -6186 709082
rect -6806 670218 -6774 670454
rect -6538 670218 -6454 670454
rect -6218 670218 -6186 670454
rect -6806 670134 -6186 670218
rect -6806 669898 -6774 670134
rect -6538 669898 -6454 670134
rect -6218 669898 -6186 670134
rect -6806 634454 -6186 669898
rect -6806 634218 -6774 634454
rect -6538 634218 -6454 634454
rect -6218 634218 -6186 634454
rect -6806 634134 -6186 634218
rect -6806 633898 -6774 634134
rect -6538 633898 -6454 634134
rect -6218 633898 -6186 634134
rect -6806 598454 -6186 633898
rect -6806 598218 -6774 598454
rect -6538 598218 -6454 598454
rect -6218 598218 -6186 598454
rect -6806 598134 -6186 598218
rect -6806 597898 -6774 598134
rect -6538 597898 -6454 598134
rect -6218 597898 -6186 598134
rect -6806 562454 -6186 597898
rect -6806 562218 -6774 562454
rect -6538 562218 -6454 562454
rect -6218 562218 -6186 562454
rect -6806 562134 -6186 562218
rect -6806 561898 -6774 562134
rect -6538 561898 -6454 562134
rect -6218 561898 -6186 562134
rect -6806 526454 -6186 561898
rect -6806 526218 -6774 526454
rect -6538 526218 -6454 526454
rect -6218 526218 -6186 526454
rect -6806 526134 -6186 526218
rect -6806 525898 -6774 526134
rect -6538 525898 -6454 526134
rect -6218 525898 -6186 526134
rect -6806 490454 -6186 525898
rect -6806 490218 -6774 490454
rect -6538 490218 -6454 490454
rect -6218 490218 -6186 490454
rect -6806 490134 -6186 490218
rect -6806 489898 -6774 490134
rect -6538 489898 -6454 490134
rect -6218 489898 -6186 490134
rect -6806 454454 -6186 489898
rect -6806 454218 -6774 454454
rect -6538 454218 -6454 454454
rect -6218 454218 -6186 454454
rect -6806 454134 -6186 454218
rect -6806 453898 -6774 454134
rect -6538 453898 -6454 454134
rect -6218 453898 -6186 454134
rect -6806 418454 -6186 453898
rect -6806 418218 -6774 418454
rect -6538 418218 -6454 418454
rect -6218 418218 -6186 418454
rect -6806 418134 -6186 418218
rect -6806 417898 -6774 418134
rect -6538 417898 -6454 418134
rect -6218 417898 -6186 418134
rect -6806 382454 -6186 417898
rect -6806 382218 -6774 382454
rect -6538 382218 -6454 382454
rect -6218 382218 -6186 382454
rect -6806 382134 -6186 382218
rect -6806 381898 -6774 382134
rect -6538 381898 -6454 382134
rect -6218 381898 -6186 382134
rect -6806 346454 -6186 381898
rect -6806 346218 -6774 346454
rect -6538 346218 -6454 346454
rect -6218 346218 -6186 346454
rect -6806 346134 -6186 346218
rect -6806 345898 -6774 346134
rect -6538 345898 -6454 346134
rect -6218 345898 -6186 346134
rect -6806 310454 -6186 345898
rect -6806 310218 -6774 310454
rect -6538 310218 -6454 310454
rect -6218 310218 -6186 310454
rect -6806 310134 -6186 310218
rect -6806 309898 -6774 310134
rect -6538 309898 -6454 310134
rect -6218 309898 -6186 310134
rect -6806 274454 -6186 309898
rect -6806 274218 -6774 274454
rect -6538 274218 -6454 274454
rect -6218 274218 -6186 274454
rect -6806 274134 -6186 274218
rect -6806 273898 -6774 274134
rect -6538 273898 -6454 274134
rect -6218 273898 -6186 274134
rect -6806 238454 -6186 273898
rect -6806 238218 -6774 238454
rect -6538 238218 -6454 238454
rect -6218 238218 -6186 238454
rect -6806 238134 -6186 238218
rect -6806 237898 -6774 238134
rect -6538 237898 -6454 238134
rect -6218 237898 -6186 238134
rect -6806 202454 -6186 237898
rect -6806 202218 -6774 202454
rect -6538 202218 -6454 202454
rect -6218 202218 -6186 202454
rect -6806 202134 -6186 202218
rect -6806 201898 -6774 202134
rect -6538 201898 -6454 202134
rect -6218 201898 -6186 202134
rect -6806 166454 -6186 201898
rect -6806 166218 -6774 166454
rect -6538 166218 -6454 166454
rect -6218 166218 -6186 166454
rect -6806 166134 -6186 166218
rect -6806 165898 -6774 166134
rect -6538 165898 -6454 166134
rect -6218 165898 -6186 166134
rect -6806 130454 -6186 165898
rect -6806 130218 -6774 130454
rect -6538 130218 -6454 130454
rect -6218 130218 -6186 130454
rect -6806 130134 -6186 130218
rect -6806 129898 -6774 130134
rect -6538 129898 -6454 130134
rect -6218 129898 -6186 130134
rect -6806 94454 -6186 129898
rect -6806 94218 -6774 94454
rect -6538 94218 -6454 94454
rect -6218 94218 -6186 94454
rect -6806 94134 -6186 94218
rect -6806 93898 -6774 94134
rect -6538 93898 -6454 94134
rect -6218 93898 -6186 94134
rect -6806 58454 -6186 93898
rect -6806 58218 -6774 58454
rect -6538 58218 -6454 58454
rect -6218 58218 -6186 58454
rect -6806 58134 -6186 58218
rect -6806 57898 -6774 58134
rect -6538 57898 -6454 58134
rect -6218 57898 -6186 58134
rect -6806 22454 -6186 57898
rect -6806 22218 -6774 22454
rect -6538 22218 -6454 22454
rect -6218 22218 -6186 22454
rect -6806 22134 -6186 22218
rect -6806 21898 -6774 22134
rect -6538 21898 -6454 22134
rect -6218 21898 -6186 22134
rect -6806 -5146 -6186 21898
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666734 -5226 708122
rect -5846 666498 -5814 666734
rect -5578 666498 -5494 666734
rect -5258 666498 -5226 666734
rect -5846 666414 -5226 666498
rect -5846 666178 -5814 666414
rect -5578 666178 -5494 666414
rect -5258 666178 -5226 666414
rect -5846 630734 -5226 666178
rect -5846 630498 -5814 630734
rect -5578 630498 -5494 630734
rect -5258 630498 -5226 630734
rect -5846 630414 -5226 630498
rect -5846 630178 -5814 630414
rect -5578 630178 -5494 630414
rect -5258 630178 -5226 630414
rect -5846 594734 -5226 630178
rect -5846 594498 -5814 594734
rect -5578 594498 -5494 594734
rect -5258 594498 -5226 594734
rect -5846 594414 -5226 594498
rect -5846 594178 -5814 594414
rect -5578 594178 -5494 594414
rect -5258 594178 -5226 594414
rect -5846 558734 -5226 594178
rect -5846 558498 -5814 558734
rect -5578 558498 -5494 558734
rect -5258 558498 -5226 558734
rect -5846 558414 -5226 558498
rect -5846 558178 -5814 558414
rect -5578 558178 -5494 558414
rect -5258 558178 -5226 558414
rect -5846 522734 -5226 558178
rect -5846 522498 -5814 522734
rect -5578 522498 -5494 522734
rect -5258 522498 -5226 522734
rect -5846 522414 -5226 522498
rect -5846 522178 -5814 522414
rect -5578 522178 -5494 522414
rect -5258 522178 -5226 522414
rect -5846 486734 -5226 522178
rect -5846 486498 -5814 486734
rect -5578 486498 -5494 486734
rect -5258 486498 -5226 486734
rect -5846 486414 -5226 486498
rect -5846 486178 -5814 486414
rect -5578 486178 -5494 486414
rect -5258 486178 -5226 486414
rect -5846 450734 -5226 486178
rect -5846 450498 -5814 450734
rect -5578 450498 -5494 450734
rect -5258 450498 -5226 450734
rect -5846 450414 -5226 450498
rect -5846 450178 -5814 450414
rect -5578 450178 -5494 450414
rect -5258 450178 -5226 450414
rect -5846 414734 -5226 450178
rect -5846 414498 -5814 414734
rect -5578 414498 -5494 414734
rect -5258 414498 -5226 414734
rect -5846 414414 -5226 414498
rect -5846 414178 -5814 414414
rect -5578 414178 -5494 414414
rect -5258 414178 -5226 414414
rect -5846 378734 -5226 414178
rect -5846 378498 -5814 378734
rect -5578 378498 -5494 378734
rect -5258 378498 -5226 378734
rect -5846 378414 -5226 378498
rect -5846 378178 -5814 378414
rect -5578 378178 -5494 378414
rect -5258 378178 -5226 378414
rect -5846 342734 -5226 378178
rect -5846 342498 -5814 342734
rect -5578 342498 -5494 342734
rect -5258 342498 -5226 342734
rect -5846 342414 -5226 342498
rect -5846 342178 -5814 342414
rect -5578 342178 -5494 342414
rect -5258 342178 -5226 342414
rect -5846 306734 -5226 342178
rect -5846 306498 -5814 306734
rect -5578 306498 -5494 306734
rect -5258 306498 -5226 306734
rect -5846 306414 -5226 306498
rect -5846 306178 -5814 306414
rect -5578 306178 -5494 306414
rect -5258 306178 -5226 306414
rect -5846 270734 -5226 306178
rect -5846 270498 -5814 270734
rect -5578 270498 -5494 270734
rect -5258 270498 -5226 270734
rect -5846 270414 -5226 270498
rect -5846 270178 -5814 270414
rect -5578 270178 -5494 270414
rect -5258 270178 -5226 270414
rect -5846 234734 -5226 270178
rect -5846 234498 -5814 234734
rect -5578 234498 -5494 234734
rect -5258 234498 -5226 234734
rect -5846 234414 -5226 234498
rect -5846 234178 -5814 234414
rect -5578 234178 -5494 234414
rect -5258 234178 -5226 234414
rect -5846 198734 -5226 234178
rect -5846 198498 -5814 198734
rect -5578 198498 -5494 198734
rect -5258 198498 -5226 198734
rect -5846 198414 -5226 198498
rect -5846 198178 -5814 198414
rect -5578 198178 -5494 198414
rect -5258 198178 -5226 198414
rect -5846 162734 -5226 198178
rect -5846 162498 -5814 162734
rect -5578 162498 -5494 162734
rect -5258 162498 -5226 162734
rect -5846 162414 -5226 162498
rect -5846 162178 -5814 162414
rect -5578 162178 -5494 162414
rect -5258 162178 -5226 162414
rect -5846 126734 -5226 162178
rect -5846 126498 -5814 126734
rect -5578 126498 -5494 126734
rect -5258 126498 -5226 126734
rect -5846 126414 -5226 126498
rect -5846 126178 -5814 126414
rect -5578 126178 -5494 126414
rect -5258 126178 -5226 126414
rect -5846 90734 -5226 126178
rect -5846 90498 -5814 90734
rect -5578 90498 -5494 90734
rect -5258 90498 -5226 90734
rect -5846 90414 -5226 90498
rect -5846 90178 -5814 90414
rect -5578 90178 -5494 90414
rect -5258 90178 -5226 90414
rect -5846 54734 -5226 90178
rect -5846 54498 -5814 54734
rect -5578 54498 -5494 54734
rect -5258 54498 -5226 54734
rect -5846 54414 -5226 54498
rect -5846 54178 -5814 54414
rect -5578 54178 -5494 54414
rect -5258 54178 -5226 54414
rect -5846 18734 -5226 54178
rect -5846 18498 -5814 18734
rect -5578 18498 -5494 18734
rect -5258 18498 -5226 18734
rect -5846 18414 -5226 18498
rect -5846 18178 -5814 18414
rect -5578 18178 -5494 18414
rect -5258 18178 -5226 18414
rect -5846 -4186 -5226 18178
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 699014 -4266 707162
rect -4886 698778 -4854 699014
rect -4618 698778 -4534 699014
rect -4298 698778 -4266 699014
rect -4886 698694 -4266 698778
rect -4886 698458 -4854 698694
rect -4618 698458 -4534 698694
rect -4298 698458 -4266 698694
rect -4886 663014 -4266 698458
rect -4886 662778 -4854 663014
rect -4618 662778 -4534 663014
rect -4298 662778 -4266 663014
rect -4886 662694 -4266 662778
rect -4886 662458 -4854 662694
rect -4618 662458 -4534 662694
rect -4298 662458 -4266 662694
rect -4886 627014 -4266 662458
rect -4886 626778 -4854 627014
rect -4618 626778 -4534 627014
rect -4298 626778 -4266 627014
rect -4886 626694 -4266 626778
rect -4886 626458 -4854 626694
rect -4618 626458 -4534 626694
rect -4298 626458 -4266 626694
rect -4886 591014 -4266 626458
rect -4886 590778 -4854 591014
rect -4618 590778 -4534 591014
rect -4298 590778 -4266 591014
rect -4886 590694 -4266 590778
rect -4886 590458 -4854 590694
rect -4618 590458 -4534 590694
rect -4298 590458 -4266 590694
rect -4886 555014 -4266 590458
rect -4886 554778 -4854 555014
rect -4618 554778 -4534 555014
rect -4298 554778 -4266 555014
rect -4886 554694 -4266 554778
rect -4886 554458 -4854 554694
rect -4618 554458 -4534 554694
rect -4298 554458 -4266 554694
rect -4886 519014 -4266 554458
rect -4886 518778 -4854 519014
rect -4618 518778 -4534 519014
rect -4298 518778 -4266 519014
rect -4886 518694 -4266 518778
rect -4886 518458 -4854 518694
rect -4618 518458 -4534 518694
rect -4298 518458 -4266 518694
rect -4886 483014 -4266 518458
rect -4886 482778 -4854 483014
rect -4618 482778 -4534 483014
rect -4298 482778 -4266 483014
rect -4886 482694 -4266 482778
rect -4886 482458 -4854 482694
rect -4618 482458 -4534 482694
rect -4298 482458 -4266 482694
rect -4886 447014 -4266 482458
rect -4886 446778 -4854 447014
rect -4618 446778 -4534 447014
rect -4298 446778 -4266 447014
rect -4886 446694 -4266 446778
rect -4886 446458 -4854 446694
rect -4618 446458 -4534 446694
rect -4298 446458 -4266 446694
rect -4886 411014 -4266 446458
rect -4886 410778 -4854 411014
rect -4618 410778 -4534 411014
rect -4298 410778 -4266 411014
rect -4886 410694 -4266 410778
rect -4886 410458 -4854 410694
rect -4618 410458 -4534 410694
rect -4298 410458 -4266 410694
rect -4886 375014 -4266 410458
rect -4886 374778 -4854 375014
rect -4618 374778 -4534 375014
rect -4298 374778 -4266 375014
rect -4886 374694 -4266 374778
rect -4886 374458 -4854 374694
rect -4618 374458 -4534 374694
rect -4298 374458 -4266 374694
rect -4886 339014 -4266 374458
rect -4886 338778 -4854 339014
rect -4618 338778 -4534 339014
rect -4298 338778 -4266 339014
rect -4886 338694 -4266 338778
rect -4886 338458 -4854 338694
rect -4618 338458 -4534 338694
rect -4298 338458 -4266 338694
rect -4886 303014 -4266 338458
rect -4886 302778 -4854 303014
rect -4618 302778 -4534 303014
rect -4298 302778 -4266 303014
rect -4886 302694 -4266 302778
rect -4886 302458 -4854 302694
rect -4618 302458 -4534 302694
rect -4298 302458 -4266 302694
rect -4886 267014 -4266 302458
rect -4886 266778 -4854 267014
rect -4618 266778 -4534 267014
rect -4298 266778 -4266 267014
rect -4886 266694 -4266 266778
rect -4886 266458 -4854 266694
rect -4618 266458 -4534 266694
rect -4298 266458 -4266 266694
rect -4886 231014 -4266 266458
rect -4886 230778 -4854 231014
rect -4618 230778 -4534 231014
rect -4298 230778 -4266 231014
rect -4886 230694 -4266 230778
rect -4886 230458 -4854 230694
rect -4618 230458 -4534 230694
rect -4298 230458 -4266 230694
rect -4886 195014 -4266 230458
rect -4886 194778 -4854 195014
rect -4618 194778 -4534 195014
rect -4298 194778 -4266 195014
rect -4886 194694 -4266 194778
rect -4886 194458 -4854 194694
rect -4618 194458 -4534 194694
rect -4298 194458 -4266 194694
rect -4886 159014 -4266 194458
rect -4886 158778 -4854 159014
rect -4618 158778 -4534 159014
rect -4298 158778 -4266 159014
rect -4886 158694 -4266 158778
rect -4886 158458 -4854 158694
rect -4618 158458 -4534 158694
rect -4298 158458 -4266 158694
rect -4886 123014 -4266 158458
rect -4886 122778 -4854 123014
rect -4618 122778 -4534 123014
rect -4298 122778 -4266 123014
rect -4886 122694 -4266 122778
rect -4886 122458 -4854 122694
rect -4618 122458 -4534 122694
rect -4298 122458 -4266 122694
rect -4886 87014 -4266 122458
rect -4886 86778 -4854 87014
rect -4618 86778 -4534 87014
rect -4298 86778 -4266 87014
rect -4886 86694 -4266 86778
rect -4886 86458 -4854 86694
rect -4618 86458 -4534 86694
rect -4298 86458 -4266 86694
rect -4886 51014 -4266 86458
rect -4886 50778 -4854 51014
rect -4618 50778 -4534 51014
rect -4298 50778 -4266 51014
rect -4886 50694 -4266 50778
rect -4886 50458 -4854 50694
rect -4618 50458 -4534 50694
rect -4298 50458 -4266 50694
rect -4886 15014 -4266 50458
rect -4886 14778 -4854 15014
rect -4618 14778 -4534 15014
rect -4298 14778 -4266 15014
rect -4886 14694 -4266 14778
rect -4886 14458 -4854 14694
rect -4618 14458 -4534 14694
rect -4298 14458 -4266 14694
rect -4886 -3226 -4266 14458
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 695294 -3306 706202
rect -3926 695058 -3894 695294
rect -3658 695058 -3574 695294
rect -3338 695058 -3306 695294
rect -3926 694974 -3306 695058
rect -3926 694738 -3894 694974
rect -3658 694738 -3574 694974
rect -3338 694738 -3306 694974
rect -3926 659294 -3306 694738
rect -3926 659058 -3894 659294
rect -3658 659058 -3574 659294
rect -3338 659058 -3306 659294
rect -3926 658974 -3306 659058
rect -3926 658738 -3894 658974
rect -3658 658738 -3574 658974
rect -3338 658738 -3306 658974
rect -3926 623294 -3306 658738
rect -3926 623058 -3894 623294
rect -3658 623058 -3574 623294
rect -3338 623058 -3306 623294
rect -3926 622974 -3306 623058
rect -3926 622738 -3894 622974
rect -3658 622738 -3574 622974
rect -3338 622738 -3306 622974
rect -3926 587294 -3306 622738
rect -3926 587058 -3894 587294
rect -3658 587058 -3574 587294
rect -3338 587058 -3306 587294
rect -3926 586974 -3306 587058
rect -3926 586738 -3894 586974
rect -3658 586738 -3574 586974
rect -3338 586738 -3306 586974
rect -3926 551294 -3306 586738
rect -3926 551058 -3894 551294
rect -3658 551058 -3574 551294
rect -3338 551058 -3306 551294
rect -3926 550974 -3306 551058
rect -3926 550738 -3894 550974
rect -3658 550738 -3574 550974
rect -3338 550738 -3306 550974
rect -3926 515294 -3306 550738
rect -3926 515058 -3894 515294
rect -3658 515058 -3574 515294
rect -3338 515058 -3306 515294
rect -3926 514974 -3306 515058
rect -3926 514738 -3894 514974
rect -3658 514738 -3574 514974
rect -3338 514738 -3306 514974
rect -3926 479294 -3306 514738
rect -3926 479058 -3894 479294
rect -3658 479058 -3574 479294
rect -3338 479058 -3306 479294
rect -3926 478974 -3306 479058
rect -3926 478738 -3894 478974
rect -3658 478738 -3574 478974
rect -3338 478738 -3306 478974
rect -3926 443294 -3306 478738
rect -3926 443058 -3894 443294
rect -3658 443058 -3574 443294
rect -3338 443058 -3306 443294
rect -3926 442974 -3306 443058
rect -3926 442738 -3894 442974
rect -3658 442738 -3574 442974
rect -3338 442738 -3306 442974
rect -3926 407294 -3306 442738
rect -3926 407058 -3894 407294
rect -3658 407058 -3574 407294
rect -3338 407058 -3306 407294
rect -3926 406974 -3306 407058
rect -3926 406738 -3894 406974
rect -3658 406738 -3574 406974
rect -3338 406738 -3306 406974
rect -3926 371294 -3306 406738
rect -3926 371058 -3894 371294
rect -3658 371058 -3574 371294
rect -3338 371058 -3306 371294
rect -3926 370974 -3306 371058
rect -3926 370738 -3894 370974
rect -3658 370738 -3574 370974
rect -3338 370738 -3306 370974
rect -3926 335294 -3306 370738
rect -3926 335058 -3894 335294
rect -3658 335058 -3574 335294
rect -3338 335058 -3306 335294
rect -3926 334974 -3306 335058
rect -3926 334738 -3894 334974
rect -3658 334738 -3574 334974
rect -3338 334738 -3306 334974
rect -3926 299294 -3306 334738
rect -3926 299058 -3894 299294
rect -3658 299058 -3574 299294
rect -3338 299058 -3306 299294
rect -3926 298974 -3306 299058
rect -3926 298738 -3894 298974
rect -3658 298738 -3574 298974
rect -3338 298738 -3306 298974
rect -3926 263294 -3306 298738
rect -3926 263058 -3894 263294
rect -3658 263058 -3574 263294
rect -3338 263058 -3306 263294
rect -3926 262974 -3306 263058
rect -3926 262738 -3894 262974
rect -3658 262738 -3574 262974
rect -3338 262738 -3306 262974
rect -3926 227294 -3306 262738
rect -3926 227058 -3894 227294
rect -3658 227058 -3574 227294
rect -3338 227058 -3306 227294
rect -3926 226974 -3306 227058
rect -3926 226738 -3894 226974
rect -3658 226738 -3574 226974
rect -3338 226738 -3306 226974
rect -3926 191294 -3306 226738
rect -3926 191058 -3894 191294
rect -3658 191058 -3574 191294
rect -3338 191058 -3306 191294
rect -3926 190974 -3306 191058
rect -3926 190738 -3894 190974
rect -3658 190738 -3574 190974
rect -3338 190738 -3306 190974
rect -3926 155294 -3306 190738
rect -3926 155058 -3894 155294
rect -3658 155058 -3574 155294
rect -3338 155058 -3306 155294
rect -3926 154974 -3306 155058
rect -3926 154738 -3894 154974
rect -3658 154738 -3574 154974
rect -3338 154738 -3306 154974
rect -3926 119294 -3306 154738
rect -3926 119058 -3894 119294
rect -3658 119058 -3574 119294
rect -3338 119058 -3306 119294
rect -3926 118974 -3306 119058
rect -3926 118738 -3894 118974
rect -3658 118738 -3574 118974
rect -3338 118738 -3306 118974
rect -3926 83294 -3306 118738
rect -3926 83058 -3894 83294
rect -3658 83058 -3574 83294
rect -3338 83058 -3306 83294
rect -3926 82974 -3306 83058
rect -3926 82738 -3894 82974
rect -3658 82738 -3574 82974
rect -3338 82738 -3306 82974
rect -3926 47294 -3306 82738
rect -3926 47058 -3894 47294
rect -3658 47058 -3574 47294
rect -3338 47058 -3306 47294
rect -3926 46974 -3306 47058
rect -3926 46738 -3894 46974
rect -3658 46738 -3574 46974
rect -3338 46738 -3306 46974
rect -3926 11294 -3306 46738
rect -3926 11058 -3894 11294
rect -3658 11058 -3574 11294
rect -3338 11058 -3306 11294
rect -3926 10974 -3306 11058
rect -3926 10738 -3894 10974
rect -3658 10738 -3574 10974
rect -3338 10738 -3306 10974
rect -3926 -2266 -3306 10738
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691574 -2346 705242
rect -2966 691338 -2934 691574
rect -2698 691338 -2614 691574
rect -2378 691338 -2346 691574
rect -2966 691254 -2346 691338
rect -2966 691018 -2934 691254
rect -2698 691018 -2614 691254
rect -2378 691018 -2346 691254
rect -2966 655574 -2346 691018
rect -2966 655338 -2934 655574
rect -2698 655338 -2614 655574
rect -2378 655338 -2346 655574
rect -2966 655254 -2346 655338
rect -2966 655018 -2934 655254
rect -2698 655018 -2614 655254
rect -2378 655018 -2346 655254
rect -2966 619574 -2346 655018
rect -2966 619338 -2934 619574
rect -2698 619338 -2614 619574
rect -2378 619338 -2346 619574
rect -2966 619254 -2346 619338
rect -2966 619018 -2934 619254
rect -2698 619018 -2614 619254
rect -2378 619018 -2346 619254
rect -2966 583574 -2346 619018
rect -2966 583338 -2934 583574
rect -2698 583338 -2614 583574
rect -2378 583338 -2346 583574
rect -2966 583254 -2346 583338
rect -2966 583018 -2934 583254
rect -2698 583018 -2614 583254
rect -2378 583018 -2346 583254
rect -2966 547574 -2346 583018
rect -2966 547338 -2934 547574
rect -2698 547338 -2614 547574
rect -2378 547338 -2346 547574
rect -2966 547254 -2346 547338
rect -2966 547018 -2934 547254
rect -2698 547018 -2614 547254
rect -2378 547018 -2346 547254
rect -2966 511574 -2346 547018
rect -2966 511338 -2934 511574
rect -2698 511338 -2614 511574
rect -2378 511338 -2346 511574
rect -2966 511254 -2346 511338
rect -2966 511018 -2934 511254
rect -2698 511018 -2614 511254
rect -2378 511018 -2346 511254
rect -2966 475574 -2346 511018
rect -2966 475338 -2934 475574
rect -2698 475338 -2614 475574
rect -2378 475338 -2346 475574
rect -2966 475254 -2346 475338
rect -2966 475018 -2934 475254
rect -2698 475018 -2614 475254
rect -2378 475018 -2346 475254
rect -2966 439574 -2346 475018
rect -2966 439338 -2934 439574
rect -2698 439338 -2614 439574
rect -2378 439338 -2346 439574
rect -2966 439254 -2346 439338
rect -2966 439018 -2934 439254
rect -2698 439018 -2614 439254
rect -2378 439018 -2346 439254
rect -2966 403574 -2346 439018
rect -2966 403338 -2934 403574
rect -2698 403338 -2614 403574
rect -2378 403338 -2346 403574
rect -2966 403254 -2346 403338
rect -2966 403018 -2934 403254
rect -2698 403018 -2614 403254
rect -2378 403018 -2346 403254
rect -2966 367574 -2346 403018
rect -2966 367338 -2934 367574
rect -2698 367338 -2614 367574
rect -2378 367338 -2346 367574
rect -2966 367254 -2346 367338
rect -2966 367018 -2934 367254
rect -2698 367018 -2614 367254
rect -2378 367018 -2346 367254
rect -2966 331574 -2346 367018
rect -2966 331338 -2934 331574
rect -2698 331338 -2614 331574
rect -2378 331338 -2346 331574
rect -2966 331254 -2346 331338
rect -2966 331018 -2934 331254
rect -2698 331018 -2614 331254
rect -2378 331018 -2346 331254
rect -2966 295574 -2346 331018
rect -2966 295338 -2934 295574
rect -2698 295338 -2614 295574
rect -2378 295338 -2346 295574
rect -2966 295254 -2346 295338
rect -2966 295018 -2934 295254
rect -2698 295018 -2614 295254
rect -2378 295018 -2346 295254
rect -2966 259574 -2346 295018
rect -2966 259338 -2934 259574
rect -2698 259338 -2614 259574
rect -2378 259338 -2346 259574
rect -2966 259254 -2346 259338
rect -2966 259018 -2934 259254
rect -2698 259018 -2614 259254
rect -2378 259018 -2346 259254
rect -2966 223574 -2346 259018
rect -2966 223338 -2934 223574
rect -2698 223338 -2614 223574
rect -2378 223338 -2346 223574
rect -2966 223254 -2346 223338
rect -2966 223018 -2934 223254
rect -2698 223018 -2614 223254
rect -2378 223018 -2346 223254
rect -2966 187574 -2346 223018
rect -2966 187338 -2934 187574
rect -2698 187338 -2614 187574
rect -2378 187338 -2346 187574
rect -2966 187254 -2346 187338
rect -2966 187018 -2934 187254
rect -2698 187018 -2614 187254
rect -2378 187018 -2346 187254
rect -2966 151574 -2346 187018
rect -2966 151338 -2934 151574
rect -2698 151338 -2614 151574
rect -2378 151338 -2346 151574
rect -2966 151254 -2346 151338
rect -2966 151018 -2934 151254
rect -2698 151018 -2614 151254
rect -2378 151018 -2346 151254
rect -2966 115574 -2346 151018
rect -2966 115338 -2934 115574
rect -2698 115338 -2614 115574
rect -2378 115338 -2346 115574
rect -2966 115254 -2346 115338
rect -2966 115018 -2934 115254
rect -2698 115018 -2614 115254
rect -2378 115018 -2346 115254
rect -2966 79574 -2346 115018
rect -2966 79338 -2934 79574
rect -2698 79338 -2614 79574
rect -2378 79338 -2346 79574
rect -2966 79254 -2346 79338
rect -2966 79018 -2934 79254
rect -2698 79018 -2614 79254
rect -2378 79018 -2346 79254
rect -2966 43574 -2346 79018
rect -2966 43338 -2934 43574
rect -2698 43338 -2614 43574
rect -2378 43338 -2346 43574
rect -2966 43254 -2346 43338
rect -2966 43018 -2934 43254
rect -2698 43018 -2614 43254
rect -2378 43018 -2346 43254
rect -2966 7574 -2346 43018
rect -2966 7338 -2934 7574
rect -2698 7338 -2614 7574
rect -2378 7338 -2346 7574
rect -2966 7254 -2346 7338
rect -2966 7018 -2934 7254
rect -2698 7018 -2614 7254
rect -2378 7018 -2346 7254
rect -2966 -1306 -2346 7018
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687854 -1386 704282
rect -2006 687618 -1974 687854
rect -1738 687618 -1654 687854
rect -1418 687618 -1386 687854
rect -2006 687534 -1386 687618
rect -2006 687298 -1974 687534
rect -1738 687298 -1654 687534
rect -1418 687298 -1386 687534
rect -2006 651854 -1386 687298
rect -2006 651618 -1974 651854
rect -1738 651618 -1654 651854
rect -1418 651618 -1386 651854
rect -2006 651534 -1386 651618
rect -2006 651298 -1974 651534
rect -1738 651298 -1654 651534
rect -1418 651298 -1386 651534
rect -2006 615854 -1386 651298
rect -2006 615618 -1974 615854
rect -1738 615618 -1654 615854
rect -1418 615618 -1386 615854
rect -2006 615534 -1386 615618
rect -2006 615298 -1974 615534
rect -1738 615298 -1654 615534
rect -1418 615298 -1386 615534
rect -2006 579854 -1386 615298
rect -2006 579618 -1974 579854
rect -1738 579618 -1654 579854
rect -1418 579618 -1386 579854
rect -2006 579534 -1386 579618
rect -2006 579298 -1974 579534
rect -1738 579298 -1654 579534
rect -1418 579298 -1386 579534
rect -2006 543854 -1386 579298
rect -2006 543618 -1974 543854
rect -1738 543618 -1654 543854
rect -1418 543618 -1386 543854
rect -2006 543534 -1386 543618
rect -2006 543298 -1974 543534
rect -1738 543298 -1654 543534
rect -1418 543298 -1386 543534
rect -2006 507854 -1386 543298
rect -2006 507618 -1974 507854
rect -1738 507618 -1654 507854
rect -1418 507618 -1386 507854
rect -2006 507534 -1386 507618
rect -2006 507298 -1974 507534
rect -1738 507298 -1654 507534
rect -1418 507298 -1386 507534
rect -2006 471854 -1386 507298
rect -2006 471618 -1974 471854
rect -1738 471618 -1654 471854
rect -1418 471618 -1386 471854
rect -2006 471534 -1386 471618
rect -2006 471298 -1974 471534
rect -1738 471298 -1654 471534
rect -1418 471298 -1386 471534
rect -2006 435854 -1386 471298
rect -2006 435618 -1974 435854
rect -1738 435618 -1654 435854
rect -1418 435618 -1386 435854
rect -2006 435534 -1386 435618
rect -2006 435298 -1974 435534
rect -1738 435298 -1654 435534
rect -1418 435298 -1386 435534
rect -2006 399854 -1386 435298
rect -2006 399618 -1974 399854
rect -1738 399618 -1654 399854
rect -1418 399618 -1386 399854
rect -2006 399534 -1386 399618
rect -2006 399298 -1974 399534
rect -1738 399298 -1654 399534
rect -1418 399298 -1386 399534
rect -2006 363854 -1386 399298
rect -2006 363618 -1974 363854
rect -1738 363618 -1654 363854
rect -1418 363618 -1386 363854
rect -2006 363534 -1386 363618
rect -2006 363298 -1974 363534
rect -1738 363298 -1654 363534
rect -1418 363298 -1386 363534
rect -2006 327854 -1386 363298
rect -2006 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 -1386 327854
rect -2006 327534 -1386 327618
rect -2006 327298 -1974 327534
rect -1738 327298 -1654 327534
rect -1418 327298 -1386 327534
rect -2006 291854 -1386 327298
rect -2006 291618 -1974 291854
rect -1738 291618 -1654 291854
rect -1418 291618 -1386 291854
rect -2006 291534 -1386 291618
rect -2006 291298 -1974 291534
rect -1738 291298 -1654 291534
rect -1418 291298 -1386 291534
rect -2006 255854 -1386 291298
rect -2006 255618 -1974 255854
rect -1738 255618 -1654 255854
rect -1418 255618 -1386 255854
rect -2006 255534 -1386 255618
rect -2006 255298 -1974 255534
rect -1738 255298 -1654 255534
rect -1418 255298 -1386 255534
rect -2006 219854 -1386 255298
rect -2006 219618 -1974 219854
rect -1738 219618 -1654 219854
rect -1418 219618 -1386 219854
rect -2006 219534 -1386 219618
rect -2006 219298 -1974 219534
rect -1738 219298 -1654 219534
rect -1418 219298 -1386 219534
rect -2006 183854 -1386 219298
rect -2006 183618 -1974 183854
rect -1738 183618 -1654 183854
rect -1418 183618 -1386 183854
rect -2006 183534 -1386 183618
rect -2006 183298 -1974 183534
rect -1738 183298 -1654 183534
rect -1418 183298 -1386 183534
rect -2006 147854 -1386 183298
rect -2006 147618 -1974 147854
rect -1738 147618 -1654 147854
rect -1418 147618 -1386 147854
rect -2006 147534 -1386 147618
rect -2006 147298 -1974 147534
rect -1738 147298 -1654 147534
rect -1418 147298 -1386 147534
rect -2006 111854 -1386 147298
rect -2006 111618 -1974 111854
rect -1738 111618 -1654 111854
rect -1418 111618 -1386 111854
rect -2006 111534 -1386 111618
rect -2006 111298 -1974 111534
rect -1738 111298 -1654 111534
rect -1418 111298 -1386 111534
rect -2006 75854 -1386 111298
rect -2006 75618 -1974 75854
rect -1738 75618 -1654 75854
rect -1418 75618 -1386 75854
rect -2006 75534 -1386 75618
rect -2006 75298 -1974 75534
rect -1738 75298 -1654 75534
rect -1418 75298 -1386 75534
rect -2006 39854 -1386 75298
rect -2006 39618 -1974 39854
rect -1738 39618 -1654 39854
rect -1418 39618 -1386 39854
rect -2006 39534 -1386 39618
rect -2006 39298 -1974 39534
rect -1738 39298 -1654 39534
rect -1418 39298 -1386 39534
rect -2006 3854 -1386 39298
rect -2006 3618 -1974 3854
rect -1738 3618 -1654 3854
rect -1418 3618 -1386 3854
rect -2006 3534 -1386 3618
rect -2006 3298 -1974 3534
rect -1738 3298 -1654 3534
rect -1418 3298 -1386 3534
rect -2006 -346 -1386 3298
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 2194 704838 2814 711590
rect 2194 704602 2226 704838
rect 2462 704602 2546 704838
rect 2782 704602 2814 704838
rect 2194 704518 2814 704602
rect 2194 704282 2226 704518
rect 2462 704282 2546 704518
rect 2782 704282 2814 704518
rect 2194 687854 2814 704282
rect 2194 687618 2226 687854
rect 2462 687618 2546 687854
rect 2782 687618 2814 687854
rect 2194 687534 2814 687618
rect 2194 687298 2226 687534
rect 2462 687298 2546 687534
rect 2782 687298 2814 687534
rect 2194 651854 2814 687298
rect 2194 651618 2226 651854
rect 2462 651618 2546 651854
rect 2782 651618 2814 651854
rect 2194 651534 2814 651618
rect 2194 651298 2226 651534
rect 2462 651298 2546 651534
rect 2782 651298 2814 651534
rect 2194 615854 2814 651298
rect 2194 615618 2226 615854
rect 2462 615618 2546 615854
rect 2782 615618 2814 615854
rect 2194 615534 2814 615618
rect 2194 615298 2226 615534
rect 2462 615298 2546 615534
rect 2782 615298 2814 615534
rect 2194 579854 2814 615298
rect 2194 579618 2226 579854
rect 2462 579618 2546 579854
rect 2782 579618 2814 579854
rect 2194 579534 2814 579618
rect 2194 579298 2226 579534
rect 2462 579298 2546 579534
rect 2782 579298 2814 579534
rect 2194 543854 2814 579298
rect 2194 543618 2226 543854
rect 2462 543618 2546 543854
rect 2782 543618 2814 543854
rect 2194 543534 2814 543618
rect 2194 543298 2226 543534
rect 2462 543298 2546 543534
rect 2782 543298 2814 543534
rect 2194 507854 2814 543298
rect 2194 507618 2226 507854
rect 2462 507618 2546 507854
rect 2782 507618 2814 507854
rect 2194 507534 2814 507618
rect 2194 507298 2226 507534
rect 2462 507298 2546 507534
rect 2782 507298 2814 507534
rect 2194 471854 2814 507298
rect 2194 471618 2226 471854
rect 2462 471618 2546 471854
rect 2782 471618 2814 471854
rect 2194 471534 2814 471618
rect 2194 471298 2226 471534
rect 2462 471298 2546 471534
rect 2782 471298 2814 471534
rect 2194 435854 2814 471298
rect 2194 435618 2226 435854
rect 2462 435618 2546 435854
rect 2782 435618 2814 435854
rect 2194 435534 2814 435618
rect 2194 435298 2226 435534
rect 2462 435298 2546 435534
rect 2782 435298 2814 435534
rect 2194 399854 2814 435298
rect 2194 399618 2226 399854
rect 2462 399618 2546 399854
rect 2782 399618 2814 399854
rect 2194 399534 2814 399618
rect 2194 399298 2226 399534
rect 2462 399298 2546 399534
rect 2782 399298 2814 399534
rect 2194 363854 2814 399298
rect 2194 363618 2226 363854
rect 2462 363618 2546 363854
rect 2782 363618 2814 363854
rect 2194 363534 2814 363618
rect 2194 363298 2226 363534
rect 2462 363298 2546 363534
rect 2782 363298 2814 363534
rect 2194 327854 2814 363298
rect 2194 327618 2226 327854
rect 2462 327618 2546 327854
rect 2782 327618 2814 327854
rect 2194 327534 2814 327618
rect 2194 327298 2226 327534
rect 2462 327298 2546 327534
rect 2782 327298 2814 327534
rect 2194 291854 2814 327298
rect 2194 291618 2226 291854
rect 2462 291618 2546 291854
rect 2782 291618 2814 291854
rect 2194 291534 2814 291618
rect 2194 291298 2226 291534
rect 2462 291298 2546 291534
rect 2782 291298 2814 291534
rect 2194 255854 2814 291298
rect 2194 255618 2226 255854
rect 2462 255618 2546 255854
rect 2782 255618 2814 255854
rect 2194 255534 2814 255618
rect 2194 255298 2226 255534
rect 2462 255298 2546 255534
rect 2782 255298 2814 255534
rect 2194 219854 2814 255298
rect 2194 219618 2226 219854
rect 2462 219618 2546 219854
rect 2782 219618 2814 219854
rect 2194 219534 2814 219618
rect 2194 219298 2226 219534
rect 2462 219298 2546 219534
rect 2782 219298 2814 219534
rect 2194 183854 2814 219298
rect 2194 183618 2226 183854
rect 2462 183618 2546 183854
rect 2782 183618 2814 183854
rect 2194 183534 2814 183618
rect 2194 183298 2226 183534
rect 2462 183298 2546 183534
rect 2782 183298 2814 183534
rect 2194 147854 2814 183298
rect 2194 147618 2226 147854
rect 2462 147618 2546 147854
rect 2782 147618 2814 147854
rect 2194 147534 2814 147618
rect 2194 147298 2226 147534
rect 2462 147298 2546 147534
rect 2782 147298 2814 147534
rect 2194 111854 2814 147298
rect 2194 111618 2226 111854
rect 2462 111618 2546 111854
rect 2782 111618 2814 111854
rect 2194 111534 2814 111618
rect 2194 111298 2226 111534
rect 2462 111298 2546 111534
rect 2782 111298 2814 111534
rect 2194 75854 2814 111298
rect 2194 75618 2226 75854
rect 2462 75618 2546 75854
rect 2782 75618 2814 75854
rect 2194 75534 2814 75618
rect 2194 75298 2226 75534
rect 2462 75298 2546 75534
rect 2782 75298 2814 75534
rect 2194 39854 2814 75298
rect 2194 39618 2226 39854
rect 2462 39618 2546 39854
rect 2782 39618 2814 39854
rect 2194 39534 2814 39618
rect 2194 39298 2226 39534
rect 2462 39298 2546 39534
rect 2782 39298 2814 39534
rect 2194 3854 2814 39298
rect 2194 3618 2226 3854
rect 2462 3618 2546 3854
rect 2782 3618 2814 3854
rect 2194 3534 2814 3618
rect 2194 3298 2226 3534
rect 2462 3298 2546 3534
rect 2782 3298 2814 3534
rect 2194 -346 2814 3298
rect 2194 -582 2226 -346
rect 2462 -582 2546 -346
rect 2782 -582 2814 -346
rect 2194 -666 2814 -582
rect 2194 -902 2226 -666
rect 2462 -902 2546 -666
rect 2782 -902 2814 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 2194 -7654 2814 -902
rect 5914 705798 6534 711590
rect 5914 705562 5946 705798
rect 6182 705562 6266 705798
rect 6502 705562 6534 705798
rect 5914 705478 6534 705562
rect 5914 705242 5946 705478
rect 6182 705242 6266 705478
rect 6502 705242 6534 705478
rect 5914 691574 6534 705242
rect 5914 691338 5946 691574
rect 6182 691338 6266 691574
rect 6502 691338 6534 691574
rect 5914 691254 6534 691338
rect 5914 691018 5946 691254
rect 6182 691018 6266 691254
rect 6502 691018 6534 691254
rect 5914 655574 6534 691018
rect 5914 655338 5946 655574
rect 6182 655338 6266 655574
rect 6502 655338 6534 655574
rect 5914 655254 6534 655338
rect 5914 655018 5946 655254
rect 6182 655018 6266 655254
rect 6502 655018 6534 655254
rect 5914 619574 6534 655018
rect 5914 619338 5946 619574
rect 6182 619338 6266 619574
rect 6502 619338 6534 619574
rect 5914 619254 6534 619338
rect 5914 619018 5946 619254
rect 6182 619018 6266 619254
rect 6502 619018 6534 619254
rect 5914 583574 6534 619018
rect 5914 583338 5946 583574
rect 6182 583338 6266 583574
rect 6502 583338 6534 583574
rect 5914 583254 6534 583338
rect 5914 583018 5946 583254
rect 6182 583018 6266 583254
rect 6502 583018 6534 583254
rect 5914 547574 6534 583018
rect 5914 547338 5946 547574
rect 6182 547338 6266 547574
rect 6502 547338 6534 547574
rect 5914 547254 6534 547338
rect 5914 547018 5946 547254
rect 6182 547018 6266 547254
rect 6502 547018 6534 547254
rect 5914 511574 6534 547018
rect 5914 511338 5946 511574
rect 6182 511338 6266 511574
rect 6502 511338 6534 511574
rect 5914 511254 6534 511338
rect 5914 511018 5946 511254
rect 6182 511018 6266 511254
rect 6502 511018 6534 511254
rect 5914 475574 6534 511018
rect 5914 475338 5946 475574
rect 6182 475338 6266 475574
rect 6502 475338 6534 475574
rect 5914 475254 6534 475338
rect 5914 475018 5946 475254
rect 6182 475018 6266 475254
rect 6502 475018 6534 475254
rect 5914 439574 6534 475018
rect 5914 439338 5946 439574
rect 6182 439338 6266 439574
rect 6502 439338 6534 439574
rect 5914 439254 6534 439338
rect 5914 439018 5946 439254
rect 6182 439018 6266 439254
rect 6502 439018 6534 439254
rect 5914 403574 6534 439018
rect 5914 403338 5946 403574
rect 6182 403338 6266 403574
rect 6502 403338 6534 403574
rect 5914 403254 6534 403338
rect 5914 403018 5946 403254
rect 6182 403018 6266 403254
rect 6502 403018 6534 403254
rect 5914 367574 6534 403018
rect 5914 367338 5946 367574
rect 6182 367338 6266 367574
rect 6502 367338 6534 367574
rect 5914 367254 6534 367338
rect 5914 367018 5946 367254
rect 6182 367018 6266 367254
rect 6502 367018 6534 367254
rect 5914 331574 6534 367018
rect 5914 331338 5946 331574
rect 6182 331338 6266 331574
rect 6502 331338 6534 331574
rect 5914 331254 6534 331338
rect 5914 331018 5946 331254
rect 6182 331018 6266 331254
rect 6502 331018 6534 331254
rect 5914 295574 6534 331018
rect 5914 295338 5946 295574
rect 6182 295338 6266 295574
rect 6502 295338 6534 295574
rect 5914 295254 6534 295338
rect 5914 295018 5946 295254
rect 6182 295018 6266 295254
rect 6502 295018 6534 295254
rect 5914 259574 6534 295018
rect 5914 259338 5946 259574
rect 6182 259338 6266 259574
rect 6502 259338 6534 259574
rect 5914 259254 6534 259338
rect 5914 259018 5946 259254
rect 6182 259018 6266 259254
rect 6502 259018 6534 259254
rect 5914 223574 6534 259018
rect 5914 223338 5946 223574
rect 6182 223338 6266 223574
rect 6502 223338 6534 223574
rect 5914 223254 6534 223338
rect 5914 223018 5946 223254
rect 6182 223018 6266 223254
rect 6502 223018 6534 223254
rect 5914 187574 6534 223018
rect 5914 187338 5946 187574
rect 6182 187338 6266 187574
rect 6502 187338 6534 187574
rect 5914 187254 6534 187338
rect 5914 187018 5946 187254
rect 6182 187018 6266 187254
rect 6502 187018 6534 187254
rect 5914 151574 6534 187018
rect 5914 151338 5946 151574
rect 6182 151338 6266 151574
rect 6502 151338 6534 151574
rect 5914 151254 6534 151338
rect 5914 151018 5946 151254
rect 6182 151018 6266 151254
rect 6502 151018 6534 151254
rect 5914 115574 6534 151018
rect 5914 115338 5946 115574
rect 6182 115338 6266 115574
rect 6502 115338 6534 115574
rect 5914 115254 6534 115338
rect 5914 115018 5946 115254
rect 6182 115018 6266 115254
rect 6502 115018 6534 115254
rect 5914 79574 6534 115018
rect 5914 79338 5946 79574
rect 6182 79338 6266 79574
rect 6502 79338 6534 79574
rect 5914 79254 6534 79338
rect 5914 79018 5946 79254
rect 6182 79018 6266 79254
rect 6502 79018 6534 79254
rect 5914 43574 6534 79018
rect 5914 43338 5946 43574
rect 6182 43338 6266 43574
rect 6502 43338 6534 43574
rect 5914 43254 6534 43338
rect 5914 43018 5946 43254
rect 6182 43018 6266 43254
rect 6502 43018 6534 43254
rect 5914 7574 6534 43018
rect 5914 7338 5946 7574
rect 6182 7338 6266 7574
rect 6502 7338 6534 7574
rect 5914 7254 6534 7338
rect 5914 7018 5946 7254
rect 6182 7018 6266 7254
rect 6502 7018 6534 7254
rect 5914 -1306 6534 7018
rect 5914 -1542 5946 -1306
rect 6182 -1542 6266 -1306
rect 6502 -1542 6534 -1306
rect 5914 -1626 6534 -1542
rect 5914 -1862 5946 -1626
rect 6182 -1862 6266 -1626
rect 6502 -1862 6534 -1626
rect 5914 -7654 6534 -1862
rect 9634 706758 10254 711590
rect 9634 706522 9666 706758
rect 9902 706522 9986 706758
rect 10222 706522 10254 706758
rect 9634 706438 10254 706522
rect 9634 706202 9666 706438
rect 9902 706202 9986 706438
rect 10222 706202 10254 706438
rect 9634 695294 10254 706202
rect 9634 695058 9666 695294
rect 9902 695058 9986 695294
rect 10222 695058 10254 695294
rect 9634 694974 10254 695058
rect 9634 694738 9666 694974
rect 9902 694738 9986 694974
rect 10222 694738 10254 694974
rect 9634 659294 10254 694738
rect 9634 659058 9666 659294
rect 9902 659058 9986 659294
rect 10222 659058 10254 659294
rect 9634 658974 10254 659058
rect 9634 658738 9666 658974
rect 9902 658738 9986 658974
rect 10222 658738 10254 658974
rect 9634 623294 10254 658738
rect 9634 623058 9666 623294
rect 9902 623058 9986 623294
rect 10222 623058 10254 623294
rect 9634 622974 10254 623058
rect 9634 622738 9666 622974
rect 9902 622738 9986 622974
rect 10222 622738 10254 622974
rect 9634 587294 10254 622738
rect 9634 587058 9666 587294
rect 9902 587058 9986 587294
rect 10222 587058 10254 587294
rect 9634 586974 10254 587058
rect 9634 586738 9666 586974
rect 9902 586738 9986 586974
rect 10222 586738 10254 586974
rect 9634 551294 10254 586738
rect 9634 551058 9666 551294
rect 9902 551058 9986 551294
rect 10222 551058 10254 551294
rect 9634 550974 10254 551058
rect 9634 550738 9666 550974
rect 9902 550738 9986 550974
rect 10222 550738 10254 550974
rect 9634 515294 10254 550738
rect 9634 515058 9666 515294
rect 9902 515058 9986 515294
rect 10222 515058 10254 515294
rect 9634 514974 10254 515058
rect 9634 514738 9666 514974
rect 9902 514738 9986 514974
rect 10222 514738 10254 514974
rect 9634 479294 10254 514738
rect 9634 479058 9666 479294
rect 9902 479058 9986 479294
rect 10222 479058 10254 479294
rect 9634 478974 10254 479058
rect 9634 478738 9666 478974
rect 9902 478738 9986 478974
rect 10222 478738 10254 478974
rect 9634 443294 10254 478738
rect 9634 443058 9666 443294
rect 9902 443058 9986 443294
rect 10222 443058 10254 443294
rect 9634 442974 10254 443058
rect 9634 442738 9666 442974
rect 9902 442738 9986 442974
rect 10222 442738 10254 442974
rect 9634 407294 10254 442738
rect 9634 407058 9666 407294
rect 9902 407058 9986 407294
rect 10222 407058 10254 407294
rect 9634 406974 10254 407058
rect 9634 406738 9666 406974
rect 9902 406738 9986 406974
rect 10222 406738 10254 406974
rect 9634 371294 10254 406738
rect 9634 371058 9666 371294
rect 9902 371058 9986 371294
rect 10222 371058 10254 371294
rect 9634 370974 10254 371058
rect 9634 370738 9666 370974
rect 9902 370738 9986 370974
rect 10222 370738 10254 370974
rect 9634 335294 10254 370738
rect 9634 335058 9666 335294
rect 9902 335058 9986 335294
rect 10222 335058 10254 335294
rect 9634 334974 10254 335058
rect 9634 334738 9666 334974
rect 9902 334738 9986 334974
rect 10222 334738 10254 334974
rect 9634 299294 10254 334738
rect 9634 299058 9666 299294
rect 9902 299058 9986 299294
rect 10222 299058 10254 299294
rect 9634 298974 10254 299058
rect 9634 298738 9666 298974
rect 9902 298738 9986 298974
rect 10222 298738 10254 298974
rect 9634 263294 10254 298738
rect 9634 263058 9666 263294
rect 9902 263058 9986 263294
rect 10222 263058 10254 263294
rect 9634 262974 10254 263058
rect 9634 262738 9666 262974
rect 9902 262738 9986 262974
rect 10222 262738 10254 262974
rect 9634 227294 10254 262738
rect 9634 227058 9666 227294
rect 9902 227058 9986 227294
rect 10222 227058 10254 227294
rect 9634 226974 10254 227058
rect 9634 226738 9666 226974
rect 9902 226738 9986 226974
rect 10222 226738 10254 226974
rect 9634 191294 10254 226738
rect 9634 191058 9666 191294
rect 9902 191058 9986 191294
rect 10222 191058 10254 191294
rect 9634 190974 10254 191058
rect 9634 190738 9666 190974
rect 9902 190738 9986 190974
rect 10222 190738 10254 190974
rect 9634 155294 10254 190738
rect 9634 155058 9666 155294
rect 9902 155058 9986 155294
rect 10222 155058 10254 155294
rect 9634 154974 10254 155058
rect 9634 154738 9666 154974
rect 9902 154738 9986 154974
rect 10222 154738 10254 154974
rect 9634 119294 10254 154738
rect 9634 119058 9666 119294
rect 9902 119058 9986 119294
rect 10222 119058 10254 119294
rect 9634 118974 10254 119058
rect 9634 118738 9666 118974
rect 9902 118738 9986 118974
rect 10222 118738 10254 118974
rect 9634 83294 10254 118738
rect 9634 83058 9666 83294
rect 9902 83058 9986 83294
rect 10222 83058 10254 83294
rect 9634 82974 10254 83058
rect 9634 82738 9666 82974
rect 9902 82738 9986 82974
rect 10222 82738 10254 82974
rect 9634 47294 10254 82738
rect 9634 47058 9666 47294
rect 9902 47058 9986 47294
rect 10222 47058 10254 47294
rect 9634 46974 10254 47058
rect 9634 46738 9666 46974
rect 9902 46738 9986 46974
rect 10222 46738 10254 46974
rect 9634 11294 10254 46738
rect 9634 11058 9666 11294
rect 9902 11058 9986 11294
rect 10222 11058 10254 11294
rect 9634 10974 10254 11058
rect 9634 10738 9666 10974
rect 9902 10738 9986 10974
rect 10222 10738 10254 10974
rect 9634 -2266 10254 10738
rect 13354 707718 13974 711590
rect 13354 707482 13386 707718
rect 13622 707482 13706 707718
rect 13942 707482 13974 707718
rect 13354 707398 13974 707482
rect 13354 707162 13386 707398
rect 13622 707162 13706 707398
rect 13942 707162 13974 707398
rect 13354 699014 13974 707162
rect 13354 698778 13386 699014
rect 13622 698778 13706 699014
rect 13942 698778 13974 699014
rect 13354 698694 13974 698778
rect 13354 698458 13386 698694
rect 13622 698458 13706 698694
rect 13942 698458 13974 698694
rect 13354 663014 13974 698458
rect 13354 662778 13386 663014
rect 13622 662778 13706 663014
rect 13942 662778 13974 663014
rect 13354 662694 13974 662778
rect 13354 662458 13386 662694
rect 13622 662458 13706 662694
rect 13942 662458 13974 662694
rect 13354 627014 13974 662458
rect 13354 626778 13386 627014
rect 13622 626778 13706 627014
rect 13942 626778 13974 627014
rect 13354 626694 13974 626778
rect 13354 626458 13386 626694
rect 13622 626458 13706 626694
rect 13942 626458 13974 626694
rect 13354 591014 13974 626458
rect 13354 590778 13386 591014
rect 13622 590778 13706 591014
rect 13942 590778 13974 591014
rect 13354 590694 13974 590778
rect 13354 590458 13386 590694
rect 13622 590458 13706 590694
rect 13942 590458 13974 590694
rect 13354 555014 13974 590458
rect 13354 554778 13386 555014
rect 13622 554778 13706 555014
rect 13942 554778 13974 555014
rect 13354 554694 13974 554778
rect 13354 554458 13386 554694
rect 13622 554458 13706 554694
rect 13942 554458 13974 554694
rect 13354 519014 13974 554458
rect 13354 518778 13386 519014
rect 13622 518778 13706 519014
rect 13942 518778 13974 519014
rect 13354 518694 13974 518778
rect 13354 518458 13386 518694
rect 13622 518458 13706 518694
rect 13942 518458 13974 518694
rect 13354 483014 13974 518458
rect 13354 482778 13386 483014
rect 13622 482778 13706 483014
rect 13942 482778 13974 483014
rect 13354 482694 13974 482778
rect 13354 482458 13386 482694
rect 13622 482458 13706 482694
rect 13942 482458 13974 482694
rect 13354 447014 13974 482458
rect 13354 446778 13386 447014
rect 13622 446778 13706 447014
rect 13942 446778 13974 447014
rect 13354 446694 13974 446778
rect 13354 446458 13386 446694
rect 13622 446458 13706 446694
rect 13942 446458 13974 446694
rect 13354 411014 13974 446458
rect 13354 410778 13386 411014
rect 13622 410778 13706 411014
rect 13942 410778 13974 411014
rect 13354 410694 13974 410778
rect 13354 410458 13386 410694
rect 13622 410458 13706 410694
rect 13942 410458 13974 410694
rect 13354 375014 13974 410458
rect 13354 374778 13386 375014
rect 13622 374778 13706 375014
rect 13942 374778 13974 375014
rect 13354 374694 13974 374778
rect 13354 374458 13386 374694
rect 13622 374458 13706 374694
rect 13942 374458 13974 374694
rect 13354 339014 13974 374458
rect 13354 338778 13386 339014
rect 13622 338778 13706 339014
rect 13942 338778 13974 339014
rect 13354 338694 13974 338778
rect 13354 338458 13386 338694
rect 13622 338458 13706 338694
rect 13942 338458 13974 338694
rect 13354 303014 13974 338458
rect 13354 302778 13386 303014
rect 13622 302778 13706 303014
rect 13942 302778 13974 303014
rect 13354 302694 13974 302778
rect 13354 302458 13386 302694
rect 13622 302458 13706 302694
rect 13942 302458 13974 302694
rect 13354 267014 13974 302458
rect 13354 266778 13386 267014
rect 13622 266778 13706 267014
rect 13942 266778 13974 267014
rect 13354 266694 13974 266778
rect 13354 266458 13386 266694
rect 13622 266458 13706 266694
rect 13942 266458 13974 266694
rect 13354 231014 13974 266458
rect 13354 230778 13386 231014
rect 13622 230778 13706 231014
rect 13942 230778 13974 231014
rect 13354 230694 13974 230778
rect 13354 230458 13386 230694
rect 13622 230458 13706 230694
rect 13942 230458 13974 230694
rect 13354 195014 13974 230458
rect 13354 194778 13386 195014
rect 13622 194778 13706 195014
rect 13942 194778 13974 195014
rect 13354 194694 13974 194778
rect 13354 194458 13386 194694
rect 13622 194458 13706 194694
rect 13942 194458 13974 194694
rect 13354 159014 13974 194458
rect 13354 158778 13386 159014
rect 13622 158778 13706 159014
rect 13942 158778 13974 159014
rect 13354 158694 13974 158778
rect 13354 158458 13386 158694
rect 13622 158458 13706 158694
rect 13942 158458 13974 158694
rect 13354 123014 13974 158458
rect 13354 122778 13386 123014
rect 13622 122778 13706 123014
rect 13942 122778 13974 123014
rect 13354 122694 13974 122778
rect 13354 122458 13386 122694
rect 13622 122458 13706 122694
rect 13942 122458 13974 122694
rect 13354 87014 13974 122458
rect 13354 86778 13386 87014
rect 13622 86778 13706 87014
rect 13942 86778 13974 87014
rect 13354 86694 13974 86778
rect 13354 86458 13386 86694
rect 13622 86458 13706 86694
rect 13942 86458 13974 86694
rect 13354 51014 13974 86458
rect 13354 50778 13386 51014
rect 13622 50778 13706 51014
rect 13942 50778 13974 51014
rect 13354 50694 13974 50778
rect 13354 50458 13386 50694
rect 13622 50458 13706 50694
rect 13942 50458 13974 50694
rect 13354 15014 13974 50458
rect 13354 14778 13386 15014
rect 13622 14778 13706 15014
rect 13942 14778 13974 15014
rect 13354 14694 13974 14778
rect 13354 14458 13386 14694
rect 13622 14458 13706 14694
rect 13942 14458 13974 14694
rect 12390 2821 12450 4302
rect 12387 2820 12453 2821
rect 12387 2756 12388 2820
rect 12452 2756 12453 2820
rect 12387 2755 12453 2756
rect 9634 -2502 9666 -2266
rect 9902 -2502 9986 -2266
rect 10222 -2502 10254 -2266
rect 9634 -2586 10254 -2502
rect 9634 -2822 9666 -2586
rect 9902 -2822 9986 -2586
rect 10222 -2822 10254 -2586
rect 9634 -7654 10254 -2822
rect 13354 -3226 13974 14458
rect 13354 -3462 13386 -3226
rect 13622 -3462 13706 -3226
rect 13942 -3462 13974 -3226
rect 13354 -3546 13974 -3462
rect 13354 -3782 13386 -3546
rect 13622 -3782 13706 -3546
rect 13942 -3782 13974 -3546
rect 13354 -7654 13974 -3782
rect 17074 708678 17694 711590
rect 17074 708442 17106 708678
rect 17342 708442 17426 708678
rect 17662 708442 17694 708678
rect 17074 708358 17694 708442
rect 17074 708122 17106 708358
rect 17342 708122 17426 708358
rect 17662 708122 17694 708358
rect 17074 666734 17694 708122
rect 17074 666498 17106 666734
rect 17342 666498 17426 666734
rect 17662 666498 17694 666734
rect 17074 666414 17694 666498
rect 17074 666178 17106 666414
rect 17342 666178 17426 666414
rect 17662 666178 17694 666414
rect 17074 630734 17694 666178
rect 17074 630498 17106 630734
rect 17342 630498 17426 630734
rect 17662 630498 17694 630734
rect 17074 630414 17694 630498
rect 17074 630178 17106 630414
rect 17342 630178 17426 630414
rect 17662 630178 17694 630414
rect 17074 594734 17694 630178
rect 17074 594498 17106 594734
rect 17342 594498 17426 594734
rect 17662 594498 17694 594734
rect 17074 594414 17694 594498
rect 17074 594178 17106 594414
rect 17342 594178 17426 594414
rect 17662 594178 17694 594414
rect 17074 558734 17694 594178
rect 17074 558498 17106 558734
rect 17342 558498 17426 558734
rect 17662 558498 17694 558734
rect 17074 558414 17694 558498
rect 17074 558178 17106 558414
rect 17342 558178 17426 558414
rect 17662 558178 17694 558414
rect 17074 522734 17694 558178
rect 17074 522498 17106 522734
rect 17342 522498 17426 522734
rect 17662 522498 17694 522734
rect 17074 522414 17694 522498
rect 17074 522178 17106 522414
rect 17342 522178 17426 522414
rect 17662 522178 17694 522414
rect 17074 486734 17694 522178
rect 17074 486498 17106 486734
rect 17342 486498 17426 486734
rect 17662 486498 17694 486734
rect 17074 486414 17694 486498
rect 17074 486178 17106 486414
rect 17342 486178 17426 486414
rect 17662 486178 17694 486414
rect 17074 450734 17694 486178
rect 17074 450498 17106 450734
rect 17342 450498 17426 450734
rect 17662 450498 17694 450734
rect 17074 450414 17694 450498
rect 17074 450178 17106 450414
rect 17342 450178 17426 450414
rect 17662 450178 17694 450414
rect 17074 414734 17694 450178
rect 17074 414498 17106 414734
rect 17342 414498 17426 414734
rect 17662 414498 17694 414734
rect 17074 414414 17694 414498
rect 17074 414178 17106 414414
rect 17342 414178 17426 414414
rect 17662 414178 17694 414414
rect 17074 378734 17694 414178
rect 17074 378498 17106 378734
rect 17342 378498 17426 378734
rect 17662 378498 17694 378734
rect 17074 378414 17694 378498
rect 17074 378178 17106 378414
rect 17342 378178 17426 378414
rect 17662 378178 17694 378414
rect 17074 342734 17694 378178
rect 17074 342498 17106 342734
rect 17342 342498 17426 342734
rect 17662 342498 17694 342734
rect 17074 342414 17694 342498
rect 17074 342178 17106 342414
rect 17342 342178 17426 342414
rect 17662 342178 17694 342414
rect 17074 306734 17694 342178
rect 17074 306498 17106 306734
rect 17342 306498 17426 306734
rect 17662 306498 17694 306734
rect 17074 306414 17694 306498
rect 17074 306178 17106 306414
rect 17342 306178 17426 306414
rect 17662 306178 17694 306414
rect 17074 270734 17694 306178
rect 17074 270498 17106 270734
rect 17342 270498 17426 270734
rect 17662 270498 17694 270734
rect 17074 270414 17694 270498
rect 17074 270178 17106 270414
rect 17342 270178 17426 270414
rect 17662 270178 17694 270414
rect 17074 234734 17694 270178
rect 17074 234498 17106 234734
rect 17342 234498 17426 234734
rect 17662 234498 17694 234734
rect 17074 234414 17694 234498
rect 17074 234178 17106 234414
rect 17342 234178 17426 234414
rect 17662 234178 17694 234414
rect 17074 198734 17694 234178
rect 17074 198498 17106 198734
rect 17342 198498 17426 198734
rect 17662 198498 17694 198734
rect 17074 198414 17694 198498
rect 17074 198178 17106 198414
rect 17342 198178 17426 198414
rect 17662 198178 17694 198414
rect 17074 162734 17694 198178
rect 17074 162498 17106 162734
rect 17342 162498 17426 162734
rect 17662 162498 17694 162734
rect 17074 162414 17694 162498
rect 17074 162178 17106 162414
rect 17342 162178 17426 162414
rect 17662 162178 17694 162414
rect 17074 126734 17694 162178
rect 17074 126498 17106 126734
rect 17342 126498 17426 126734
rect 17662 126498 17694 126734
rect 17074 126414 17694 126498
rect 17074 126178 17106 126414
rect 17342 126178 17426 126414
rect 17662 126178 17694 126414
rect 17074 90734 17694 126178
rect 17074 90498 17106 90734
rect 17342 90498 17426 90734
rect 17662 90498 17694 90734
rect 17074 90414 17694 90498
rect 17074 90178 17106 90414
rect 17342 90178 17426 90414
rect 17662 90178 17694 90414
rect 17074 54734 17694 90178
rect 17074 54498 17106 54734
rect 17342 54498 17426 54734
rect 17662 54498 17694 54734
rect 17074 54414 17694 54498
rect 17074 54178 17106 54414
rect 17342 54178 17426 54414
rect 17662 54178 17694 54414
rect 17074 18734 17694 54178
rect 17074 18498 17106 18734
rect 17342 18498 17426 18734
rect 17662 18498 17694 18734
rect 17074 18414 17694 18498
rect 17074 18178 17106 18414
rect 17342 18178 17426 18414
rect 17662 18178 17694 18414
rect 17074 -4186 17694 18178
rect 17074 -4422 17106 -4186
rect 17342 -4422 17426 -4186
rect 17662 -4422 17694 -4186
rect 17074 -4506 17694 -4422
rect 17074 -4742 17106 -4506
rect 17342 -4742 17426 -4506
rect 17662 -4742 17694 -4506
rect 17074 -7654 17694 -4742
rect 20794 709638 21414 711590
rect 20794 709402 20826 709638
rect 21062 709402 21146 709638
rect 21382 709402 21414 709638
rect 20794 709318 21414 709402
rect 20794 709082 20826 709318
rect 21062 709082 21146 709318
rect 21382 709082 21414 709318
rect 20794 670454 21414 709082
rect 20794 670218 20826 670454
rect 21062 670218 21146 670454
rect 21382 670218 21414 670454
rect 20794 670134 21414 670218
rect 20794 669898 20826 670134
rect 21062 669898 21146 670134
rect 21382 669898 21414 670134
rect 20794 634454 21414 669898
rect 20794 634218 20826 634454
rect 21062 634218 21146 634454
rect 21382 634218 21414 634454
rect 20794 634134 21414 634218
rect 20794 633898 20826 634134
rect 21062 633898 21146 634134
rect 21382 633898 21414 634134
rect 20794 598454 21414 633898
rect 20794 598218 20826 598454
rect 21062 598218 21146 598454
rect 21382 598218 21414 598454
rect 20794 598134 21414 598218
rect 20794 597898 20826 598134
rect 21062 597898 21146 598134
rect 21382 597898 21414 598134
rect 20794 562454 21414 597898
rect 20794 562218 20826 562454
rect 21062 562218 21146 562454
rect 21382 562218 21414 562454
rect 20794 562134 21414 562218
rect 20794 561898 20826 562134
rect 21062 561898 21146 562134
rect 21382 561898 21414 562134
rect 20794 526454 21414 561898
rect 20794 526218 20826 526454
rect 21062 526218 21146 526454
rect 21382 526218 21414 526454
rect 20794 526134 21414 526218
rect 20794 525898 20826 526134
rect 21062 525898 21146 526134
rect 21382 525898 21414 526134
rect 20794 490454 21414 525898
rect 20794 490218 20826 490454
rect 21062 490218 21146 490454
rect 21382 490218 21414 490454
rect 20794 490134 21414 490218
rect 20794 489898 20826 490134
rect 21062 489898 21146 490134
rect 21382 489898 21414 490134
rect 20794 454454 21414 489898
rect 20794 454218 20826 454454
rect 21062 454218 21146 454454
rect 21382 454218 21414 454454
rect 20794 454134 21414 454218
rect 20794 453898 20826 454134
rect 21062 453898 21146 454134
rect 21382 453898 21414 454134
rect 20794 418454 21414 453898
rect 20794 418218 20826 418454
rect 21062 418218 21146 418454
rect 21382 418218 21414 418454
rect 20794 418134 21414 418218
rect 20794 417898 20826 418134
rect 21062 417898 21146 418134
rect 21382 417898 21414 418134
rect 20794 382454 21414 417898
rect 20794 382218 20826 382454
rect 21062 382218 21146 382454
rect 21382 382218 21414 382454
rect 20794 382134 21414 382218
rect 20794 381898 20826 382134
rect 21062 381898 21146 382134
rect 21382 381898 21414 382134
rect 20794 346454 21414 381898
rect 20794 346218 20826 346454
rect 21062 346218 21146 346454
rect 21382 346218 21414 346454
rect 20794 346134 21414 346218
rect 20794 345898 20826 346134
rect 21062 345898 21146 346134
rect 21382 345898 21414 346134
rect 20794 310454 21414 345898
rect 20794 310218 20826 310454
rect 21062 310218 21146 310454
rect 21382 310218 21414 310454
rect 20794 310134 21414 310218
rect 20794 309898 20826 310134
rect 21062 309898 21146 310134
rect 21382 309898 21414 310134
rect 20794 274454 21414 309898
rect 20794 274218 20826 274454
rect 21062 274218 21146 274454
rect 21382 274218 21414 274454
rect 20794 274134 21414 274218
rect 20794 273898 20826 274134
rect 21062 273898 21146 274134
rect 21382 273898 21414 274134
rect 20794 238454 21414 273898
rect 20794 238218 20826 238454
rect 21062 238218 21146 238454
rect 21382 238218 21414 238454
rect 20794 238134 21414 238218
rect 20794 237898 20826 238134
rect 21062 237898 21146 238134
rect 21382 237898 21414 238134
rect 20794 202454 21414 237898
rect 20794 202218 20826 202454
rect 21062 202218 21146 202454
rect 21382 202218 21414 202454
rect 20794 202134 21414 202218
rect 20794 201898 20826 202134
rect 21062 201898 21146 202134
rect 21382 201898 21414 202134
rect 20794 166454 21414 201898
rect 20794 166218 20826 166454
rect 21062 166218 21146 166454
rect 21382 166218 21414 166454
rect 20794 166134 21414 166218
rect 20794 165898 20826 166134
rect 21062 165898 21146 166134
rect 21382 165898 21414 166134
rect 20794 130454 21414 165898
rect 20794 130218 20826 130454
rect 21062 130218 21146 130454
rect 21382 130218 21414 130454
rect 20794 130134 21414 130218
rect 20794 129898 20826 130134
rect 21062 129898 21146 130134
rect 21382 129898 21414 130134
rect 20794 94454 21414 129898
rect 20794 94218 20826 94454
rect 21062 94218 21146 94454
rect 21382 94218 21414 94454
rect 20794 94134 21414 94218
rect 20794 93898 20826 94134
rect 21062 93898 21146 94134
rect 21382 93898 21414 94134
rect 20794 58454 21414 93898
rect 20794 58218 20826 58454
rect 21062 58218 21146 58454
rect 21382 58218 21414 58454
rect 20794 58134 21414 58218
rect 20794 57898 20826 58134
rect 21062 57898 21146 58134
rect 21382 57898 21414 58134
rect 20794 22454 21414 57898
rect 20794 22218 20826 22454
rect 21062 22218 21146 22454
rect 21382 22218 21414 22454
rect 20794 22134 21414 22218
rect 20794 21898 20826 22134
rect 21062 21898 21146 22134
rect 21382 21898 21414 22134
rect 20794 -5146 21414 21898
rect 20794 -5382 20826 -5146
rect 21062 -5382 21146 -5146
rect 21382 -5382 21414 -5146
rect 20794 -5466 21414 -5382
rect 20794 -5702 20826 -5466
rect 21062 -5702 21146 -5466
rect 21382 -5702 21414 -5466
rect 20794 -7654 21414 -5702
rect 24514 710598 25134 711590
rect 24514 710362 24546 710598
rect 24782 710362 24866 710598
rect 25102 710362 25134 710598
rect 24514 710278 25134 710362
rect 24514 710042 24546 710278
rect 24782 710042 24866 710278
rect 25102 710042 25134 710278
rect 24514 674174 25134 710042
rect 24514 673938 24546 674174
rect 24782 673938 24866 674174
rect 25102 673938 25134 674174
rect 24514 673854 25134 673938
rect 24514 673618 24546 673854
rect 24782 673618 24866 673854
rect 25102 673618 25134 673854
rect 24514 638174 25134 673618
rect 24514 637938 24546 638174
rect 24782 637938 24866 638174
rect 25102 637938 25134 638174
rect 24514 637854 25134 637938
rect 24514 637618 24546 637854
rect 24782 637618 24866 637854
rect 25102 637618 25134 637854
rect 24514 602174 25134 637618
rect 24514 601938 24546 602174
rect 24782 601938 24866 602174
rect 25102 601938 25134 602174
rect 24514 601854 25134 601938
rect 24514 601618 24546 601854
rect 24782 601618 24866 601854
rect 25102 601618 25134 601854
rect 24514 566174 25134 601618
rect 24514 565938 24546 566174
rect 24782 565938 24866 566174
rect 25102 565938 25134 566174
rect 24514 565854 25134 565938
rect 24514 565618 24546 565854
rect 24782 565618 24866 565854
rect 25102 565618 25134 565854
rect 24514 530174 25134 565618
rect 24514 529938 24546 530174
rect 24782 529938 24866 530174
rect 25102 529938 25134 530174
rect 24514 529854 25134 529938
rect 24514 529618 24546 529854
rect 24782 529618 24866 529854
rect 25102 529618 25134 529854
rect 24514 494174 25134 529618
rect 24514 493938 24546 494174
rect 24782 493938 24866 494174
rect 25102 493938 25134 494174
rect 24514 493854 25134 493938
rect 24514 493618 24546 493854
rect 24782 493618 24866 493854
rect 25102 493618 25134 493854
rect 24514 458174 25134 493618
rect 24514 457938 24546 458174
rect 24782 457938 24866 458174
rect 25102 457938 25134 458174
rect 24514 457854 25134 457938
rect 24514 457618 24546 457854
rect 24782 457618 24866 457854
rect 25102 457618 25134 457854
rect 24514 422174 25134 457618
rect 24514 421938 24546 422174
rect 24782 421938 24866 422174
rect 25102 421938 25134 422174
rect 24514 421854 25134 421938
rect 24514 421618 24546 421854
rect 24782 421618 24866 421854
rect 25102 421618 25134 421854
rect 24514 386174 25134 421618
rect 24514 385938 24546 386174
rect 24782 385938 24866 386174
rect 25102 385938 25134 386174
rect 24514 385854 25134 385938
rect 24514 385618 24546 385854
rect 24782 385618 24866 385854
rect 25102 385618 25134 385854
rect 24514 350174 25134 385618
rect 24514 349938 24546 350174
rect 24782 349938 24866 350174
rect 25102 349938 25134 350174
rect 24514 349854 25134 349938
rect 24514 349618 24546 349854
rect 24782 349618 24866 349854
rect 25102 349618 25134 349854
rect 24514 314174 25134 349618
rect 24514 313938 24546 314174
rect 24782 313938 24866 314174
rect 25102 313938 25134 314174
rect 24514 313854 25134 313938
rect 24514 313618 24546 313854
rect 24782 313618 24866 313854
rect 25102 313618 25134 313854
rect 24514 278174 25134 313618
rect 24514 277938 24546 278174
rect 24782 277938 24866 278174
rect 25102 277938 25134 278174
rect 24514 277854 25134 277938
rect 24514 277618 24546 277854
rect 24782 277618 24866 277854
rect 25102 277618 25134 277854
rect 24514 242174 25134 277618
rect 24514 241938 24546 242174
rect 24782 241938 24866 242174
rect 25102 241938 25134 242174
rect 24514 241854 25134 241938
rect 24514 241618 24546 241854
rect 24782 241618 24866 241854
rect 25102 241618 25134 241854
rect 24514 206174 25134 241618
rect 24514 205938 24546 206174
rect 24782 205938 24866 206174
rect 25102 205938 25134 206174
rect 24514 205854 25134 205938
rect 24514 205618 24546 205854
rect 24782 205618 24866 205854
rect 25102 205618 25134 205854
rect 24514 170174 25134 205618
rect 24514 169938 24546 170174
rect 24782 169938 24866 170174
rect 25102 169938 25134 170174
rect 24514 169854 25134 169938
rect 24514 169618 24546 169854
rect 24782 169618 24866 169854
rect 25102 169618 25134 169854
rect 24514 134174 25134 169618
rect 24514 133938 24546 134174
rect 24782 133938 24866 134174
rect 25102 133938 25134 134174
rect 24514 133854 25134 133938
rect 24514 133618 24546 133854
rect 24782 133618 24866 133854
rect 25102 133618 25134 133854
rect 24514 98174 25134 133618
rect 24514 97938 24546 98174
rect 24782 97938 24866 98174
rect 25102 97938 25134 98174
rect 24514 97854 25134 97938
rect 24514 97618 24546 97854
rect 24782 97618 24866 97854
rect 25102 97618 25134 97854
rect 24514 62174 25134 97618
rect 24514 61938 24546 62174
rect 24782 61938 24866 62174
rect 25102 61938 25134 62174
rect 24514 61854 25134 61938
rect 24514 61618 24546 61854
rect 24782 61618 24866 61854
rect 25102 61618 25134 61854
rect 24514 26174 25134 61618
rect 24514 25938 24546 26174
rect 24782 25938 24866 26174
rect 25102 25938 25134 26174
rect 24514 25854 25134 25938
rect 24514 25618 24546 25854
rect 24782 25618 24866 25854
rect 25102 25618 25134 25854
rect 24514 -6106 25134 25618
rect 28234 711558 28854 711590
rect 28234 711322 28266 711558
rect 28502 711322 28586 711558
rect 28822 711322 28854 711558
rect 28234 711238 28854 711322
rect 28234 711002 28266 711238
rect 28502 711002 28586 711238
rect 28822 711002 28854 711238
rect 28234 677894 28854 711002
rect 28234 677658 28266 677894
rect 28502 677658 28586 677894
rect 28822 677658 28854 677894
rect 28234 677574 28854 677658
rect 28234 677338 28266 677574
rect 28502 677338 28586 677574
rect 28822 677338 28854 677574
rect 28234 641894 28854 677338
rect 28234 641658 28266 641894
rect 28502 641658 28586 641894
rect 28822 641658 28854 641894
rect 28234 641574 28854 641658
rect 28234 641338 28266 641574
rect 28502 641338 28586 641574
rect 28822 641338 28854 641574
rect 28234 605894 28854 641338
rect 28234 605658 28266 605894
rect 28502 605658 28586 605894
rect 28822 605658 28854 605894
rect 28234 605574 28854 605658
rect 28234 605338 28266 605574
rect 28502 605338 28586 605574
rect 28822 605338 28854 605574
rect 28234 569894 28854 605338
rect 28234 569658 28266 569894
rect 28502 569658 28586 569894
rect 28822 569658 28854 569894
rect 28234 569574 28854 569658
rect 28234 569338 28266 569574
rect 28502 569338 28586 569574
rect 28822 569338 28854 569574
rect 28234 533894 28854 569338
rect 28234 533658 28266 533894
rect 28502 533658 28586 533894
rect 28822 533658 28854 533894
rect 28234 533574 28854 533658
rect 28234 533338 28266 533574
rect 28502 533338 28586 533574
rect 28822 533338 28854 533574
rect 28234 497894 28854 533338
rect 28234 497658 28266 497894
rect 28502 497658 28586 497894
rect 28822 497658 28854 497894
rect 28234 497574 28854 497658
rect 28234 497338 28266 497574
rect 28502 497338 28586 497574
rect 28822 497338 28854 497574
rect 28234 461894 28854 497338
rect 28234 461658 28266 461894
rect 28502 461658 28586 461894
rect 28822 461658 28854 461894
rect 28234 461574 28854 461658
rect 28234 461338 28266 461574
rect 28502 461338 28586 461574
rect 28822 461338 28854 461574
rect 28234 425894 28854 461338
rect 28234 425658 28266 425894
rect 28502 425658 28586 425894
rect 28822 425658 28854 425894
rect 28234 425574 28854 425658
rect 28234 425338 28266 425574
rect 28502 425338 28586 425574
rect 28822 425338 28854 425574
rect 28234 389894 28854 425338
rect 28234 389658 28266 389894
rect 28502 389658 28586 389894
rect 28822 389658 28854 389894
rect 28234 389574 28854 389658
rect 28234 389338 28266 389574
rect 28502 389338 28586 389574
rect 28822 389338 28854 389574
rect 28234 353894 28854 389338
rect 28234 353658 28266 353894
rect 28502 353658 28586 353894
rect 28822 353658 28854 353894
rect 28234 353574 28854 353658
rect 28234 353338 28266 353574
rect 28502 353338 28586 353574
rect 28822 353338 28854 353574
rect 28234 317894 28854 353338
rect 28234 317658 28266 317894
rect 28502 317658 28586 317894
rect 28822 317658 28854 317894
rect 28234 317574 28854 317658
rect 28234 317338 28266 317574
rect 28502 317338 28586 317574
rect 28822 317338 28854 317574
rect 28234 281894 28854 317338
rect 28234 281658 28266 281894
rect 28502 281658 28586 281894
rect 28822 281658 28854 281894
rect 28234 281574 28854 281658
rect 28234 281338 28266 281574
rect 28502 281338 28586 281574
rect 28822 281338 28854 281574
rect 28234 245894 28854 281338
rect 28234 245658 28266 245894
rect 28502 245658 28586 245894
rect 28822 245658 28854 245894
rect 28234 245574 28854 245658
rect 28234 245338 28266 245574
rect 28502 245338 28586 245574
rect 28822 245338 28854 245574
rect 28234 209894 28854 245338
rect 28234 209658 28266 209894
rect 28502 209658 28586 209894
rect 28822 209658 28854 209894
rect 28234 209574 28854 209658
rect 28234 209338 28266 209574
rect 28502 209338 28586 209574
rect 28822 209338 28854 209574
rect 28234 173894 28854 209338
rect 28234 173658 28266 173894
rect 28502 173658 28586 173894
rect 28822 173658 28854 173894
rect 28234 173574 28854 173658
rect 28234 173338 28266 173574
rect 28502 173338 28586 173574
rect 28822 173338 28854 173574
rect 28234 137894 28854 173338
rect 28234 137658 28266 137894
rect 28502 137658 28586 137894
rect 28822 137658 28854 137894
rect 28234 137574 28854 137658
rect 28234 137338 28266 137574
rect 28502 137338 28586 137574
rect 28822 137338 28854 137574
rect 28234 101894 28854 137338
rect 28234 101658 28266 101894
rect 28502 101658 28586 101894
rect 28822 101658 28854 101894
rect 28234 101574 28854 101658
rect 28234 101338 28266 101574
rect 28502 101338 28586 101574
rect 28822 101338 28854 101574
rect 28234 65894 28854 101338
rect 28234 65658 28266 65894
rect 28502 65658 28586 65894
rect 28822 65658 28854 65894
rect 28234 65574 28854 65658
rect 28234 65338 28266 65574
rect 28502 65338 28586 65574
rect 28822 65338 28854 65574
rect 28234 29894 28854 65338
rect 28234 29658 28266 29894
rect 28502 29658 28586 29894
rect 28822 29658 28854 29894
rect 28234 29574 28854 29658
rect 28234 29338 28266 29574
rect 28502 29338 28586 29574
rect 28822 29338 28854 29574
rect 27846 3501 27906 9742
rect 27843 3500 27909 3501
rect 27843 3436 27844 3500
rect 27908 3436 27909 3500
rect 27843 3435 27909 3436
rect 24514 -6342 24546 -6106
rect 24782 -6342 24866 -6106
rect 25102 -6342 25134 -6106
rect 24514 -6426 25134 -6342
rect 24514 -6662 24546 -6426
rect 24782 -6662 24866 -6426
rect 25102 -6662 25134 -6426
rect 24514 -7654 25134 -6662
rect 28234 -7066 28854 29338
rect 28234 -7302 28266 -7066
rect 28502 -7302 28586 -7066
rect 28822 -7302 28854 -7066
rect 28234 -7386 28854 -7302
rect 28234 -7622 28266 -7386
rect 28502 -7622 28586 -7386
rect 28822 -7622 28854 -7386
rect 28234 -7654 28854 -7622
rect 38194 704838 38814 711590
rect 38194 704602 38226 704838
rect 38462 704602 38546 704838
rect 38782 704602 38814 704838
rect 38194 704518 38814 704602
rect 38194 704282 38226 704518
rect 38462 704282 38546 704518
rect 38782 704282 38814 704518
rect 38194 687854 38814 704282
rect 38194 687618 38226 687854
rect 38462 687618 38546 687854
rect 38782 687618 38814 687854
rect 38194 687534 38814 687618
rect 38194 687298 38226 687534
rect 38462 687298 38546 687534
rect 38782 687298 38814 687534
rect 38194 651854 38814 687298
rect 38194 651618 38226 651854
rect 38462 651618 38546 651854
rect 38782 651618 38814 651854
rect 38194 651534 38814 651618
rect 38194 651298 38226 651534
rect 38462 651298 38546 651534
rect 38782 651298 38814 651534
rect 38194 615854 38814 651298
rect 38194 615618 38226 615854
rect 38462 615618 38546 615854
rect 38782 615618 38814 615854
rect 38194 615534 38814 615618
rect 38194 615298 38226 615534
rect 38462 615298 38546 615534
rect 38782 615298 38814 615534
rect 38194 579854 38814 615298
rect 38194 579618 38226 579854
rect 38462 579618 38546 579854
rect 38782 579618 38814 579854
rect 38194 579534 38814 579618
rect 38194 579298 38226 579534
rect 38462 579298 38546 579534
rect 38782 579298 38814 579534
rect 38194 543854 38814 579298
rect 38194 543618 38226 543854
rect 38462 543618 38546 543854
rect 38782 543618 38814 543854
rect 38194 543534 38814 543618
rect 38194 543298 38226 543534
rect 38462 543298 38546 543534
rect 38782 543298 38814 543534
rect 38194 507854 38814 543298
rect 38194 507618 38226 507854
rect 38462 507618 38546 507854
rect 38782 507618 38814 507854
rect 38194 507534 38814 507618
rect 38194 507298 38226 507534
rect 38462 507298 38546 507534
rect 38782 507298 38814 507534
rect 38194 471854 38814 507298
rect 38194 471618 38226 471854
rect 38462 471618 38546 471854
rect 38782 471618 38814 471854
rect 38194 471534 38814 471618
rect 38194 471298 38226 471534
rect 38462 471298 38546 471534
rect 38782 471298 38814 471534
rect 38194 435854 38814 471298
rect 38194 435618 38226 435854
rect 38462 435618 38546 435854
rect 38782 435618 38814 435854
rect 38194 435534 38814 435618
rect 38194 435298 38226 435534
rect 38462 435298 38546 435534
rect 38782 435298 38814 435534
rect 38194 399854 38814 435298
rect 38194 399618 38226 399854
rect 38462 399618 38546 399854
rect 38782 399618 38814 399854
rect 38194 399534 38814 399618
rect 38194 399298 38226 399534
rect 38462 399298 38546 399534
rect 38782 399298 38814 399534
rect 38194 363854 38814 399298
rect 38194 363618 38226 363854
rect 38462 363618 38546 363854
rect 38782 363618 38814 363854
rect 38194 363534 38814 363618
rect 38194 363298 38226 363534
rect 38462 363298 38546 363534
rect 38782 363298 38814 363534
rect 38194 327854 38814 363298
rect 38194 327618 38226 327854
rect 38462 327618 38546 327854
rect 38782 327618 38814 327854
rect 38194 327534 38814 327618
rect 38194 327298 38226 327534
rect 38462 327298 38546 327534
rect 38782 327298 38814 327534
rect 38194 291854 38814 327298
rect 38194 291618 38226 291854
rect 38462 291618 38546 291854
rect 38782 291618 38814 291854
rect 38194 291534 38814 291618
rect 38194 291298 38226 291534
rect 38462 291298 38546 291534
rect 38782 291298 38814 291534
rect 38194 255854 38814 291298
rect 38194 255618 38226 255854
rect 38462 255618 38546 255854
rect 38782 255618 38814 255854
rect 38194 255534 38814 255618
rect 38194 255298 38226 255534
rect 38462 255298 38546 255534
rect 38782 255298 38814 255534
rect 38194 219854 38814 255298
rect 38194 219618 38226 219854
rect 38462 219618 38546 219854
rect 38782 219618 38814 219854
rect 38194 219534 38814 219618
rect 38194 219298 38226 219534
rect 38462 219298 38546 219534
rect 38782 219298 38814 219534
rect 38194 183854 38814 219298
rect 38194 183618 38226 183854
rect 38462 183618 38546 183854
rect 38782 183618 38814 183854
rect 38194 183534 38814 183618
rect 38194 183298 38226 183534
rect 38462 183298 38546 183534
rect 38782 183298 38814 183534
rect 38194 147854 38814 183298
rect 38194 147618 38226 147854
rect 38462 147618 38546 147854
rect 38782 147618 38814 147854
rect 38194 147534 38814 147618
rect 38194 147298 38226 147534
rect 38462 147298 38546 147534
rect 38782 147298 38814 147534
rect 38194 111854 38814 147298
rect 38194 111618 38226 111854
rect 38462 111618 38546 111854
rect 38782 111618 38814 111854
rect 38194 111534 38814 111618
rect 38194 111298 38226 111534
rect 38462 111298 38546 111534
rect 38782 111298 38814 111534
rect 38194 75854 38814 111298
rect 38194 75618 38226 75854
rect 38462 75618 38546 75854
rect 38782 75618 38814 75854
rect 38194 75534 38814 75618
rect 38194 75298 38226 75534
rect 38462 75298 38546 75534
rect 38782 75298 38814 75534
rect 38194 39854 38814 75298
rect 38194 39618 38226 39854
rect 38462 39618 38546 39854
rect 38782 39618 38814 39854
rect 38194 39534 38814 39618
rect 38194 39298 38226 39534
rect 38462 39298 38546 39534
rect 38782 39298 38814 39534
rect 38194 3854 38814 39298
rect 38194 3618 38226 3854
rect 38462 3618 38546 3854
rect 38782 3618 38814 3854
rect 38194 3534 38814 3618
rect 38194 3298 38226 3534
rect 38462 3298 38546 3534
rect 38782 3298 38814 3534
rect 38194 -346 38814 3298
rect 38194 -582 38226 -346
rect 38462 -582 38546 -346
rect 38782 -582 38814 -346
rect 38194 -666 38814 -582
rect 38194 -902 38226 -666
rect 38462 -902 38546 -666
rect 38782 -902 38814 -666
rect 38194 -7654 38814 -902
rect 41914 705798 42534 711590
rect 41914 705562 41946 705798
rect 42182 705562 42266 705798
rect 42502 705562 42534 705798
rect 41914 705478 42534 705562
rect 41914 705242 41946 705478
rect 42182 705242 42266 705478
rect 42502 705242 42534 705478
rect 41914 691574 42534 705242
rect 41914 691338 41946 691574
rect 42182 691338 42266 691574
rect 42502 691338 42534 691574
rect 41914 691254 42534 691338
rect 41914 691018 41946 691254
rect 42182 691018 42266 691254
rect 42502 691018 42534 691254
rect 41914 655574 42534 691018
rect 41914 655338 41946 655574
rect 42182 655338 42266 655574
rect 42502 655338 42534 655574
rect 41914 655254 42534 655338
rect 41914 655018 41946 655254
rect 42182 655018 42266 655254
rect 42502 655018 42534 655254
rect 41914 619574 42534 655018
rect 41914 619338 41946 619574
rect 42182 619338 42266 619574
rect 42502 619338 42534 619574
rect 41914 619254 42534 619338
rect 41914 619018 41946 619254
rect 42182 619018 42266 619254
rect 42502 619018 42534 619254
rect 41914 583574 42534 619018
rect 41914 583338 41946 583574
rect 42182 583338 42266 583574
rect 42502 583338 42534 583574
rect 41914 583254 42534 583338
rect 41914 583018 41946 583254
rect 42182 583018 42266 583254
rect 42502 583018 42534 583254
rect 41914 547574 42534 583018
rect 41914 547338 41946 547574
rect 42182 547338 42266 547574
rect 42502 547338 42534 547574
rect 41914 547254 42534 547338
rect 41914 547018 41946 547254
rect 42182 547018 42266 547254
rect 42502 547018 42534 547254
rect 41914 511574 42534 547018
rect 41914 511338 41946 511574
rect 42182 511338 42266 511574
rect 42502 511338 42534 511574
rect 41914 511254 42534 511338
rect 41914 511018 41946 511254
rect 42182 511018 42266 511254
rect 42502 511018 42534 511254
rect 41914 475574 42534 511018
rect 41914 475338 41946 475574
rect 42182 475338 42266 475574
rect 42502 475338 42534 475574
rect 41914 475254 42534 475338
rect 41914 475018 41946 475254
rect 42182 475018 42266 475254
rect 42502 475018 42534 475254
rect 41914 439574 42534 475018
rect 41914 439338 41946 439574
rect 42182 439338 42266 439574
rect 42502 439338 42534 439574
rect 41914 439254 42534 439338
rect 41914 439018 41946 439254
rect 42182 439018 42266 439254
rect 42502 439018 42534 439254
rect 41914 403574 42534 439018
rect 41914 403338 41946 403574
rect 42182 403338 42266 403574
rect 42502 403338 42534 403574
rect 41914 403254 42534 403338
rect 41914 403018 41946 403254
rect 42182 403018 42266 403254
rect 42502 403018 42534 403254
rect 41914 367574 42534 403018
rect 41914 367338 41946 367574
rect 42182 367338 42266 367574
rect 42502 367338 42534 367574
rect 41914 367254 42534 367338
rect 41914 367018 41946 367254
rect 42182 367018 42266 367254
rect 42502 367018 42534 367254
rect 41914 331574 42534 367018
rect 41914 331338 41946 331574
rect 42182 331338 42266 331574
rect 42502 331338 42534 331574
rect 41914 331254 42534 331338
rect 41914 331018 41946 331254
rect 42182 331018 42266 331254
rect 42502 331018 42534 331254
rect 41914 295574 42534 331018
rect 41914 295338 41946 295574
rect 42182 295338 42266 295574
rect 42502 295338 42534 295574
rect 41914 295254 42534 295338
rect 41914 295018 41946 295254
rect 42182 295018 42266 295254
rect 42502 295018 42534 295254
rect 41914 259574 42534 295018
rect 41914 259338 41946 259574
rect 42182 259338 42266 259574
rect 42502 259338 42534 259574
rect 41914 259254 42534 259338
rect 41914 259018 41946 259254
rect 42182 259018 42266 259254
rect 42502 259018 42534 259254
rect 41914 223574 42534 259018
rect 41914 223338 41946 223574
rect 42182 223338 42266 223574
rect 42502 223338 42534 223574
rect 41914 223254 42534 223338
rect 41914 223018 41946 223254
rect 42182 223018 42266 223254
rect 42502 223018 42534 223254
rect 41914 187574 42534 223018
rect 41914 187338 41946 187574
rect 42182 187338 42266 187574
rect 42502 187338 42534 187574
rect 41914 187254 42534 187338
rect 41914 187018 41946 187254
rect 42182 187018 42266 187254
rect 42502 187018 42534 187254
rect 41914 151574 42534 187018
rect 41914 151338 41946 151574
rect 42182 151338 42266 151574
rect 42502 151338 42534 151574
rect 41914 151254 42534 151338
rect 41914 151018 41946 151254
rect 42182 151018 42266 151254
rect 42502 151018 42534 151254
rect 41914 115574 42534 151018
rect 41914 115338 41946 115574
rect 42182 115338 42266 115574
rect 42502 115338 42534 115574
rect 41914 115254 42534 115338
rect 41914 115018 41946 115254
rect 42182 115018 42266 115254
rect 42502 115018 42534 115254
rect 41914 79574 42534 115018
rect 41914 79338 41946 79574
rect 42182 79338 42266 79574
rect 42502 79338 42534 79574
rect 41914 79254 42534 79338
rect 41914 79018 41946 79254
rect 42182 79018 42266 79254
rect 42502 79018 42534 79254
rect 41914 43574 42534 79018
rect 41914 43338 41946 43574
rect 42182 43338 42266 43574
rect 42502 43338 42534 43574
rect 41914 43254 42534 43338
rect 41914 43018 41946 43254
rect 42182 43018 42266 43254
rect 42502 43018 42534 43254
rect 41914 7574 42534 43018
rect 41914 7338 41946 7574
rect 42182 7338 42266 7574
rect 42502 7338 42534 7574
rect 41914 7254 42534 7338
rect 41914 7018 41946 7254
rect 42182 7018 42266 7254
rect 42502 7018 42534 7254
rect 41914 -1306 42534 7018
rect 45634 706758 46254 711590
rect 45634 706522 45666 706758
rect 45902 706522 45986 706758
rect 46222 706522 46254 706758
rect 45634 706438 46254 706522
rect 45634 706202 45666 706438
rect 45902 706202 45986 706438
rect 46222 706202 46254 706438
rect 45634 695294 46254 706202
rect 45634 695058 45666 695294
rect 45902 695058 45986 695294
rect 46222 695058 46254 695294
rect 45634 694974 46254 695058
rect 45634 694738 45666 694974
rect 45902 694738 45986 694974
rect 46222 694738 46254 694974
rect 45634 659294 46254 694738
rect 45634 659058 45666 659294
rect 45902 659058 45986 659294
rect 46222 659058 46254 659294
rect 45634 658974 46254 659058
rect 45634 658738 45666 658974
rect 45902 658738 45986 658974
rect 46222 658738 46254 658974
rect 45634 623294 46254 658738
rect 45634 623058 45666 623294
rect 45902 623058 45986 623294
rect 46222 623058 46254 623294
rect 45634 622974 46254 623058
rect 45634 622738 45666 622974
rect 45902 622738 45986 622974
rect 46222 622738 46254 622974
rect 45634 587294 46254 622738
rect 45634 587058 45666 587294
rect 45902 587058 45986 587294
rect 46222 587058 46254 587294
rect 45634 586974 46254 587058
rect 45634 586738 45666 586974
rect 45902 586738 45986 586974
rect 46222 586738 46254 586974
rect 45634 551294 46254 586738
rect 45634 551058 45666 551294
rect 45902 551058 45986 551294
rect 46222 551058 46254 551294
rect 45634 550974 46254 551058
rect 45634 550738 45666 550974
rect 45902 550738 45986 550974
rect 46222 550738 46254 550974
rect 45634 515294 46254 550738
rect 45634 515058 45666 515294
rect 45902 515058 45986 515294
rect 46222 515058 46254 515294
rect 45634 514974 46254 515058
rect 45634 514738 45666 514974
rect 45902 514738 45986 514974
rect 46222 514738 46254 514974
rect 45634 479294 46254 514738
rect 45634 479058 45666 479294
rect 45902 479058 45986 479294
rect 46222 479058 46254 479294
rect 45634 478974 46254 479058
rect 45634 478738 45666 478974
rect 45902 478738 45986 478974
rect 46222 478738 46254 478974
rect 45634 443294 46254 478738
rect 45634 443058 45666 443294
rect 45902 443058 45986 443294
rect 46222 443058 46254 443294
rect 45634 442974 46254 443058
rect 45634 442738 45666 442974
rect 45902 442738 45986 442974
rect 46222 442738 46254 442974
rect 45634 407294 46254 442738
rect 45634 407058 45666 407294
rect 45902 407058 45986 407294
rect 46222 407058 46254 407294
rect 45634 406974 46254 407058
rect 45634 406738 45666 406974
rect 45902 406738 45986 406974
rect 46222 406738 46254 406974
rect 45634 371294 46254 406738
rect 45634 371058 45666 371294
rect 45902 371058 45986 371294
rect 46222 371058 46254 371294
rect 45634 370974 46254 371058
rect 45634 370738 45666 370974
rect 45902 370738 45986 370974
rect 46222 370738 46254 370974
rect 45634 335294 46254 370738
rect 45634 335058 45666 335294
rect 45902 335058 45986 335294
rect 46222 335058 46254 335294
rect 45634 334974 46254 335058
rect 45634 334738 45666 334974
rect 45902 334738 45986 334974
rect 46222 334738 46254 334974
rect 45634 299294 46254 334738
rect 45634 299058 45666 299294
rect 45902 299058 45986 299294
rect 46222 299058 46254 299294
rect 45634 298974 46254 299058
rect 45634 298738 45666 298974
rect 45902 298738 45986 298974
rect 46222 298738 46254 298974
rect 45634 263294 46254 298738
rect 45634 263058 45666 263294
rect 45902 263058 45986 263294
rect 46222 263058 46254 263294
rect 45634 262974 46254 263058
rect 45634 262738 45666 262974
rect 45902 262738 45986 262974
rect 46222 262738 46254 262974
rect 45634 227294 46254 262738
rect 45634 227058 45666 227294
rect 45902 227058 45986 227294
rect 46222 227058 46254 227294
rect 45634 226974 46254 227058
rect 45634 226738 45666 226974
rect 45902 226738 45986 226974
rect 46222 226738 46254 226974
rect 45634 191294 46254 226738
rect 45634 191058 45666 191294
rect 45902 191058 45986 191294
rect 46222 191058 46254 191294
rect 45634 190974 46254 191058
rect 45634 190738 45666 190974
rect 45902 190738 45986 190974
rect 46222 190738 46254 190974
rect 45634 155294 46254 190738
rect 45634 155058 45666 155294
rect 45902 155058 45986 155294
rect 46222 155058 46254 155294
rect 45634 154974 46254 155058
rect 45634 154738 45666 154974
rect 45902 154738 45986 154974
rect 46222 154738 46254 154974
rect 45634 119294 46254 154738
rect 45634 119058 45666 119294
rect 45902 119058 45986 119294
rect 46222 119058 46254 119294
rect 45634 118974 46254 119058
rect 45634 118738 45666 118974
rect 45902 118738 45986 118974
rect 46222 118738 46254 118974
rect 45634 83294 46254 118738
rect 45634 83058 45666 83294
rect 45902 83058 45986 83294
rect 46222 83058 46254 83294
rect 45634 82974 46254 83058
rect 45634 82738 45666 82974
rect 45902 82738 45986 82974
rect 46222 82738 46254 82974
rect 45634 47294 46254 82738
rect 45634 47058 45666 47294
rect 45902 47058 45986 47294
rect 46222 47058 46254 47294
rect 45634 46974 46254 47058
rect 45634 46738 45666 46974
rect 45902 46738 45986 46974
rect 46222 46738 46254 46974
rect 45634 11294 46254 46738
rect 45634 11058 45666 11294
rect 45902 11058 45986 11294
rect 46222 11058 46254 11294
rect 45634 10974 46254 11058
rect 45634 10738 45666 10974
rect 45902 10738 45986 10974
rect 46222 10738 46254 10974
rect 44038 3229 44098 5662
rect 44035 3228 44101 3229
rect 44035 3164 44036 3228
rect 44100 3164 44101 3228
rect 44035 3163 44101 3164
rect 41914 -1542 41946 -1306
rect 42182 -1542 42266 -1306
rect 42502 -1542 42534 -1306
rect 41914 -1626 42534 -1542
rect 41914 -1862 41946 -1626
rect 42182 -1862 42266 -1626
rect 42502 -1862 42534 -1626
rect 41914 -7654 42534 -1862
rect 45634 -2266 46254 10738
rect 45634 -2502 45666 -2266
rect 45902 -2502 45986 -2266
rect 46222 -2502 46254 -2266
rect 45634 -2586 46254 -2502
rect 45634 -2822 45666 -2586
rect 45902 -2822 45986 -2586
rect 46222 -2822 46254 -2586
rect 45634 -7654 46254 -2822
rect 49354 707718 49974 711590
rect 49354 707482 49386 707718
rect 49622 707482 49706 707718
rect 49942 707482 49974 707718
rect 49354 707398 49974 707482
rect 49354 707162 49386 707398
rect 49622 707162 49706 707398
rect 49942 707162 49974 707398
rect 49354 699014 49974 707162
rect 49354 698778 49386 699014
rect 49622 698778 49706 699014
rect 49942 698778 49974 699014
rect 49354 698694 49974 698778
rect 49354 698458 49386 698694
rect 49622 698458 49706 698694
rect 49942 698458 49974 698694
rect 49354 663014 49974 698458
rect 49354 662778 49386 663014
rect 49622 662778 49706 663014
rect 49942 662778 49974 663014
rect 49354 662694 49974 662778
rect 49354 662458 49386 662694
rect 49622 662458 49706 662694
rect 49942 662458 49974 662694
rect 49354 627014 49974 662458
rect 49354 626778 49386 627014
rect 49622 626778 49706 627014
rect 49942 626778 49974 627014
rect 49354 626694 49974 626778
rect 49354 626458 49386 626694
rect 49622 626458 49706 626694
rect 49942 626458 49974 626694
rect 49354 591014 49974 626458
rect 49354 590778 49386 591014
rect 49622 590778 49706 591014
rect 49942 590778 49974 591014
rect 49354 590694 49974 590778
rect 49354 590458 49386 590694
rect 49622 590458 49706 590694
rect 49942 590458 49974 590694
rect 49354 555014 49974 590458
rect 49354 554778 49386 555014
rect 49622 554778 49706 555014
rect 49942 554778 49974 555014
rect 49354 554694 49974 554778
rect 49354 554458 49386 554694
rect 49622 554458 49706 554694
rect 49942 554458 49974 554694
rect 49354 519014 49974 554458
rect 49354 518778 49386 519014
rect 49622 518778 49706 519014
rect 49942 518778 49974 519014
rect 49354 518694 49974 518778
rect 49354 518458 49386 518694
rect 49622 518458 49706 518694
rect 49942 518458 49974 518694
rect 49354 483014 49974 518458
rect 49354 482778 49386 483014
rect 49622 482778 49706 483014
rect 49942 482778 49974 483014
rect 49354 482694 49974 482778
rect 49354 482458 49386 482694
rect 49622 482458 49706 482694
rect 49942 482458 49974 482694
rect 49354 447014 49974 482458
rect 49354 446778 49386 447014
rect 49622 446778 49706 447014
rect 49942 446778 49974 447014
rect 49354 446694 49974 446778
rect 49354 446458 49386 446694
rect 49622 446458 49706 446694
rect 49942 446458 49974 446694
rect 49354 411014 49974 446458
rect 49354 410778 49386 411014
rect 49622 410778 49706 411014
rect 49942 410778 49974 411014
rect 49354 410694 49974 410778
rect 49354 410458 49386 410694
rect 49622 410458 49706 410694
rect 49942 410458 49974 410694
rect 49354 375014 49974 410458
rect 49354 374778 49386 375014
rect 49622 374778 49706 375014
rect 49942 374778 49974 375014
rect 49354 374694 49974 374778
rect 49354 374458 49386 374694
rect 49622 374458 49706 374694
rect 49942 374458 49974 374694
rect 49354 339014 49974 374458
rect 49354 338778 49386 339014
rect 49622 338778 49706 339014
rect 49942 338778 49974 339014
rect 49354 338694 49974 338778
rect 49354 338458 49386 338694
rect 49622 338458 49706 338694
rect 49942 338458 49974 338694
rect 49354 303014 49974 338458
rect 49354 302778 49386 303014
rect 49622 302778 49706 303014
rect 49942 302778 49974 303014
rect 49354 302694 49974 302778
rect 49354 302458 49386 302694
rect 49622 302458 49706 302694
rect 49942 302458 49974 302694
rect 49354 267014 49974 302458
rect 49354 266778 49386 267014
rect 49622 266778 49706 267014
rect 49942 266778 49974 267014
rect 49354 266694 49974 266778
rect 49354 266458 49386 266694
rect 49622 266458 49706 266694
rect 49942 266458 49974 266694
rect 49354 231014 49974 266458
rect 49354 230778 49386 231014
rect 49622 230778 49706 231014
rect 49942 230778 49974 231014
rect 49354 230694 49974 230778
rect 49354 230458 49386 230694
rect 49622 230458 49706 230694
rect 49942 230458 49974 230694
rect 49354 195014 49974 230458
rect 49354 194778 49386 195014
rect 49622 194778 49706 195014
rect 49942 194778 49974 195014
rect 49354 194694 49974 194778
rect 49354 194458 49386 194694
rect 49622 194458 49706 194694
rect 49942 194458 49974 194694
rect 49354 159014 49974 194458
rect 49354 158778 49386 159014
rect 49622 158778 49706 159014
rect 49942 158778 49974 159014
rect 49354 158694 49974 158778
rect 49354 158458 49386 158694
rect 49622 158458 49706 158694
rect 49942 158458 49974 158694
rect 49354 123014 49974 158458
rect 49354 122778 49386 123014
rect 49622 122778 49706 123014
rect 49942 122778 49974 123014
rect 49354 122694 49974 122778
rect 49354 122458 49386 122694
rect 49622 122458 49706 122694
rect 49942 122458 49974 122694
rect 49354 87014 49974 122458
rect 49354 86778 49386 87014
rect 49622 86778 49706 87014
rect 49942 86778 49974 87014
rect 49354 86694 49974 86778
rect 49354 86458 49386 86694
rect 49622 86458 49706 86694
rect 49942 86458 49974 86694
rect 49354 51014 49974 86458
rect 49354 50778 49386 51014
rect 49622 50778 49706 51014
rect 49942 50778 49974 51014
rect 49354 50694 49974 50778
rect 49354 50458 49386 50694
rect 49622 50458 49706 50694
rect 49942 50458 49974 50694
rect 49354 15014 49974 50458
rect 49354 14778 49386 15014
rect 49622 14778 49706 15014
rect 49942 14778 49974 15014
rect 49354 14694 49974 14778
rect 49354 14458 49386 14694
rect 49622 14458 49706 14694
rect 49942 14458 49974 14694
rect 49354 -3226 49974 14458
rect 49354 -3462 49386 -3226
rect 49622 -3462 49706 -3226
rect 49942 -3462 49974 -3226
rect 49354 -3546 49974 -3462
rect 49354 -3782 49386 -3546
rect 49622 -3782 49706 -3546
rect 49942 -3782 49974 -3546
rect 49354 -7654 49974 -3782
rect 53074 708678 53694 711590
rect 53074 708442 53106 708678
rect 53342 708442 53426 708678
rect 53662 708442 53694 708678
rect 53074 708358 53694 708442
rect 53074 708122 53106 708358
rect 53342 708122 53426 708358
rect 53662 708122 53694 708358
rect 53074 666734 53694 708122
rect 53074 666498 53106 666734
rect 53342 666498 53426 666734
rect 53662 666498 53694 666734
rect 53074 666414 53694 666498
rect 53074 666178 53106 666414
rect 53342 666178 53426 666414
rect 53662 666178 53694 666414
rect 53074 630734 53694 666178
rect 53074 630498 53106 630734
rect 53342 630498 53426 630734
rect 53662 630498 53694 630734
rect 53074 630414 53694 630498
rect 53074 630178 53106 630414
rect 53342 630178 53426 630414
rect 53662 630178 53694 630414
rect 53074 594734 53694 630178
rect 53074 594498 53106 594734
rect 53342 594498 53426 594734
rect 53662 594498 53694 594734
rect 53074 594414 53694 594498
rect 53074 594178 53106 594414
rect 53342 594178 53426 594414
rect 53662 594178 53694 594414
rect 53074 558734 53694 594178
rect 53074 558498 53106 558734
rect 53342 558498 53426 558734
rect 53662 558498 53694 558734
rect 53074 558414 53694 558498
rect 53074 558178 53106 558414
rect 53342 558178 53426 558414
rect 53662 558178 53694 558414
rect 53074 522734 53694 558178
rect 53074 522498 53106 522734
rect 53342 522498 53426 522734
rect 53662 522498 53694 522734
rect 53074 522414 53694 522498
rect 53074 522178 53106 522414
rect 53342 522178 53426 522414
rect 53662 522178 53694 522414
rect 53074 486734 53694 522178
rect 53074 486498 53106 486734
rect 53342 486498 53426 486734
rect 53662 486498 53694 486734
rect 53074 486414 53694 486498
rect 53074 486178 53106 486414
rect 53342 486178 53426 486414
rect 53662 486178 53694 486414
rect 53074 450734 53694 486178
rect 53074 450498 53106 450734
rect 53342 450498 53426 450734
rect 53662 450498 53694 450734
rect 53074 450414 53694 450498
rect 53074 450178 53106 450414
rect 53342 450178 53426 450414
rect 53662 450178 53694 450414
rect 53074 414734 53694 450178
rect 53074 414498 53106 414734
rect 53342 414498 53426 414734
rect 53662 414498 53694 414734
rect 53074 414414 53694 414498
rect 53074 414178 53106 414414
rect 53342 414178 53426 414414
rect 53662 414178 53694 414414
rect 53074 378734 53694 414178
rect 53074 378498 53106 378734
rect 53342 378498 53426 378734
rect 53662 378498 53694 378734
rect 53074 378414 53694 378498
rect 53074 378178 53106 378414
rect 53342 378178 53426 378414
rect 53662 378178 53694 378414
rect 53074 342734 53694 378178
rect 53074 342498 53106 342734
rect 53342 342498 53426 342734
rect 53662 342498 53694 342734
rect 53074 342414 53694 342498
rect 53074 342178 53106 342414
rect 53342 342178 53426 342414
rect 53662 342178 53694 342414
rect 53074 306734 53694 342178
rect 53074 306498 53106 306734
rect 53342 306498 53426 306734
rect 53662 306498 53694 306734
rect 53074 306414 53694 306498
rect 53074 306178 53106 306414
rect 53342 306178 53426 306414
rect 53662 306178 53694 306414
rect 53074 270734 53694 306178
rect 53074 270498 53106 270734
rect 53342 270498 53426 270734
rect 53662 270498 53694 270734
rect 53074 270414 53694 270498
rect 53074 270178 53106 270414
rect 53342 270178 53426 270414
rect 53662 270178 53694 270414
rect 53074 234734 53694 270178
rect 53074 234498 53106 234734
rect 53342 234498 53426 234734
rect 53662 234498 53694 234734
rect 53074 234414 53694 234498
rect 53074 234178 53106 234414
rect 53342 234178 53426 234414
rect 53662 234178 53694 234414
rect 53074 198734 53694 234178
rect 53074 198498 53106 198734
rect 53342 198498 53426 198734
rect 53662 198498 53694 198734
rect 53074 198414 53694 198498
rect 53074 198178 53106 198414
rect 53342 198178 53426 198414
rect 53662 198178 53694 198414
rect 53074 162734 53694 198178
rect 53074 162498 53106 162734
rect 53342 162498 53426 162734
rect 53662 162498 53694 162734
rect 53074 162414 53694 162498
rect 53074 162178 53106 162414
rect 53342 162178 53426 162414
rect 53662 162178 53694 162414
rect 53074 126734 53694 162178
rect 53074 126498 53106 126734
rect 53342 126498 53426 126734
rect 53662 126498 53694 126734
rect 53074 126414 53694 126498
rect 53074 126178 53106 126414
rect 53342 126178 53426 126414
rect 53662 126178 53694 126414
rect 53074 90734 53694 126178
rect 53074 90498 53106 90734
rect 53342 90498 53426 90734
rect 53662 90498 53694 90734
rect 53074 90414 53694 90498
rect 53074 90178 53106 90414
rect 53342 90178 53426 90414
rect 53662 90178 53694 90414
rect 53074 54734 53694 90178
rect 53074 54498 53106 54734
rect 53342 54498 53426 54734
rect 53662 54498 53694 54734
rect 53074 54414 53694 54498
rect 53074 54178 53106 54414
rect 53342 54178 53426 54414
rect 53662 54178 53694 54414
rect 53074 18734 53694 54178
rect 53074 18498 53106 18734
rect 53342 18498 53426 18734
rect 53662 18498 53694 18734
rect 53074 18414 53694 18498
rect 53074 18178 53106 18414
rect 53342 18178 53426 18414
rect 53662 18178 53694 18414
rect 53074 -4186 53694 18178
rect 53074 -4422 53106 -4186
rect 53342 -4422 53426 -4186
rect 53662 -4422 53694 -4186
rect 53074 -4506 53694 -4422
rect 53074 -4742 53106 -4506
rect 53342 -4742 53426 -4506
rect 53662 -4742 53694 -4506
rect 53074 -7654 53694 -4742
rect 56794 709638 57414 711590
rect 56794 709402 56826 709638
rect 57062 709402 57146 709638
rect 57382 709402 57414 709638
rect 56794 709318 57414 709402
rect 56794 709082 56826 709318
rect 57062 709082 57146 709318
rect 57382 709082 57414 709318
rect 56794 670454 57414 709082
rect 56794 670218 56826 670454
rect 57062 670218 57146 670454
rect 57382 670218 57414 670454
rect 56794 670134 57414 670218
rect 56794 669898 56826 670134
rect 57062 669898 57146 670134
rect 57382 669898 57414 670134
rect 56794 634454 57414 669898
rect 56794 634218 56826 634454
rect 57062 634218 57146 634454
rect 57382 634218 57414 634454
rect 56794 634134 57414 634218
rect 56794 633898 56826 634134
rect 57062 633898 57146 634134
rect 57382 633898 57414 634134
rect 56794 598454 57414 633898
rect 56794 598218 56826 598454
rect 57062 598218 57146 598454
rect 57382 598218 57414 598454
rect 56794 598134 57414 598218
rect 56794 597898 56826 598134
rect 57062 597898 57146 598134
rect 57382 597898 57414 598134
rect 56794 562454 57414 597898
rect 56794 562218 56826 562454
rect 57062 562218 57146 562454
rect 57382 562218 57414 562454
rect 56794 562134 57414 562218
rect 56794 561898 56826 562134
rect 57062 561898 57146 562134
rect 57382 561898 57414 562134
rect 56794 526454 57414 561898
rect 56794 526218 56826 526454
rect 57062 526218 57146 526454
rect 57382 526218 57414 526454
rect 56794 526134 57414 526218
rect 56794 525898 56826 526134
rect 57062 525898 57146 526134
rect 57382 525898 57414 526134
rect 56794 490454 57414 525898
rect 56794 490218 56826 490454
rect 57062 490218 57146 490454
rect 57382 490218 57414 490454
rect 56794 490134 57414 490218
rect 56794 489898 56826 490134
rect 57062 489898 57146 490134
rect 57382 489898 57414 490134
rect 56794 454454 57414 489898
rect 56794 454218 56826 454454
rect 57062 454218 57146 454454
rect 57382 454218 57414 454454
rect 56794 454134 57414 454218
rect 56794 453898 56826 454134
rect 57062 453898 57146 454134
rect 57382 453898 57414 454134
rect 56794 418454 57414 453898
rect 56794 418218 56826 418454
rect 57062 418218 57146 418454
rect 57382 418218 57414 418454
rect 56794 418134 57414 418218
rect 56794 417898 56826 418134
rect 57062 417898 57146 418134
rect 57382 417898 57414 418134
rect 56794 382454 57414 417898
rect 56794 382218 56826 382454
rect 57062 382218 57146 382454
rect 57382 382218 57414 382454
rect 56794 382134 57414 382218
rect 56794 381898 56826 382134
rect 57062 381898 57146 382134
rect 57382 381898 57414 382134
rect 56794 346454 57414 381898
rect 56794 346218 56826 346454
rect 57062 346218 57146 346454
rect 57382 346218 57414 346454
rect 56794 346134 57414 346218
rect 56794 345898 56826 346134
rect 57062 345898 57146 346134
rect 57382 345898 57414 346134
rect 56794 310454 57414 345898
rect 56794 310218 56826 310454
rect 57062 310218 57146 310454
rect 57382 310218 57414 310454
rect 56794 310134 57414 310218
rect 56794 309898 56826 310134
rect 57062 309898 57146 310134
rect 57382 309898 57414 310134
rect 56794 274454 57414 309898
rect 56794 274218 56826 274454
rect 57062 274218 57146 274454
rect 57382 274218 57414 274454
rect 56794 274134 57414 274218
rect 56794 273898 56826 274134
rect 57062 273898 57146 274134
rect 57382 273898 57414 274134
rect 56794 238454 57414 273898
rect 56794 238218 56826 238454
rect 57062 238218 57146 238454
rect 57382 238218 57414 238454
rect 56794 238134 57414 238218
rect 56794 237898 56826 238134
rect 57062 237898 57146 238134
rect 57382 237898 57414 238134
rect 56794 202454 57414 237898
rect 56794 202218 56826 202454
rect 57062 202218 57146 202454
rect 57382 202218 57414 202454
rect 56794 202134 57414 202218
rect 56794 201898 56826 202134
rect 57062 201898 57146 202134
rect 57382 201898 57414 202134
rect 56794 166454 57414 201898
rect 56794 166218 56826 166454
rect 57062 166218 57146 166454
rect 57382 166218 57414 166454
rect 56794 166134 57414 166218
rect 56794 165898 56826 166134
rect 57062 165898 57146 166134
rect 57382 165898 57414 166134
rect 56794 130454 57414 165898
rect 56794 130218 56826 130454
rect 57062 130218 57146 130454
rect 57382 130218 57414 130454
rect 56794 130134 57414 130218
rect 56794 129898 56826 130134
rect 57062 129898 57146 130134
rect 57382 129898 57414 130134
rect 56794 94454 57414 129898
rect 56794 94218 56826 94454
rect 57062 94218 57146 94454
rect 57382 94218 57414 94454
rect 56794 94134 57414 94218
rect 56794 93898 56826 94134
rect 57062 93898 57146 94134
rect 57382 93898 57414 94134
rect 56794 58454 57414 93898
rect 56794 58218 56826 58454
rect 57062 58218 57146 58454
rect 57382 58218 57414 58454
rect 56794 58134 57414 58218
rect 56794 57898 56826 58134
rect 57062 57898 57146 58134
rect 57382 57898 57414 58134
rect 56794 22454 57414 57898
rect 56794 22218 56826 22454
rect 57062 22218 57146 22454
rect 57382 22218 57414 22454
rect 56794 22134 57414 22218
rect 56794 21898 56826 22134
rect 57062 21898 57146 22134
rect 57382 21898 57414 22134
rect 56794 -5146 57414 21898
rect 60514 710598 61134 711590
rect 60514 710362 60546 710598
rect 60782 710362 60866 710598
rect 61102 710362 61134 710598
rect 60514 710278 61134 710362
rect 60514 710042 60546 710278
rect 60782 710042 60866 710278
rect 61102 710042 61134 710278
rect 60514 674174 61134 710042
rect 60514 673938 60546 674174
rect 60782 673938 60866 674174
rect 61102 673938 61134 674174
rect 60514 673854 61134 673938
rect 60514 673618 60546 673854
rect 60782 673618 60866 673854
rect 61102 673618 61134 673854
rect 60514 638174 61134 673618
rect 60514 637938 60546 638174
rect 60782 637938 60866 638174
rect 61102 637938 61134 638174
rect 60514 637854 61134 637938
rect 60514 637618 60546 637854
rect 60782 637618 60866 637854
rect 61102 637618 61134 637854
rect 60514 602174 61134 637618
rect 60514 601938 60546 602174
rect 60782 601938 60866 602174
rect 61102 601938 61134 602174
rect 60514 601854 61134 601938
rect 60514 601618 60546 601854
rect 60782 601618 60866 601854
rect 61102 601618 61134 601854
rect 60514 566174 61134 601618
rect 60514 565938 60546 566174
rect 60782 565938 60866 566174
rect 61102 565938 61134 566174
rect 60514 565854 61134 565938
rect 60514 565618 60546 565854
rect 60782 565618 60866 565854
rect 61102 565618 61134 565854
rect 60514 530174 61134 565618
rect 60514 529938 60546 530174
rect 60782 529938 60866 530174
rect 61102 529938 61134 530174
rect 60514 529854 61134 529938
rect 60514 529618 60546 529854
rect 60782 529618 60866 529854
rect 61102 529618 61134 529854
rect 60514 494174 61134 529618
rect 60514 493938 60546 494174
rect 60782 493938 60866 494174
rect 61102 493938 61134 494174
rect 60514 493854 61134 493938
rect 60514 493618 60546 493854
rect 60782 493618 60866 493854
rect 61102 493618 61134 493854
rect 60514 458174 61134 493618
rect 60514 457938 60546 458174
rect 60782 457938 60866 458174
rect 61102 457938 61134 458174
rect 60514 457854 61134 457938
rect 60514 457618 60546 457854
rect 60782 457618 60866 457854
rect 61102 457618 61134 457854
rect 60514 422174 61134 457618
rect 60514 421938 60546 422174
rect 60782 421938 60866 422174
rect 61102 421938 61134 422174
rect 60514 421854 61134 421938
rect 60514 421618 60546 421854
rect 60782 421618 60866 421854
rect 61102 421618 61134 421854
rect 60514 386174 61134 421618
rect 60514 385938 60546 386174
rect 60782 385938 60866 386174
rect 61102 385938 61134 386174
rect 60514 385854 61134 385938
rect 60514 385618 60546 385854
rect 60782 385618 60866 385854
rect 61102 385618 61134 385854
rect 60514 350174 61134 385618
rect 60514 349938 60546 350174
rect 60782 349938 60866 350174
rect 61102 349938 61134 350174
rect 60514 349854 61134 349938
rect 60514 349618 60546 349854
rect 60782 349618 60866 349854
rect 61102 349618 61134 349854
rect 60514 314174 61134 349618
rect 60514 313938 60546 314174
rect 60782 313938 60866 314174
rect 61102 313938 61134 314174
rect 60514 313854 61134 313938
rect 60514 313618 60546 313854
rect 60782 313618 60866 313854
rect 61102 313618 61134 313854
rect 60514 278174 61134 313618
rect 60514 277938 60546 278174
rect 60782 277938 60866 278174
rect 61102 277938 61134 278174
rect 60514 277854 61134 277938
rect 60514 277618 60546 277854
rect 60782 277618 60866 277854
rect 61102 277618 61134 277854
rect 60514 242174 61134 277618
rect 60514 241938 60546 242174
rect 60782 241938 60866 242174
rect 61102 241938 61134 242174
rect 60514 241854 61134 241938
rect 60514 241618 60546 241854
rect 60782 241618 60866 241854
rect 61102 241618 61134 241854
rect 60514 206174 61134 241618
rect 60514 205938 60546 206174
rect 60782 205938 60866 206174
rect 61102 205938 61134 206174
rect 60514 205854 61134 205938
rect 60514 205618 60546 205854
rect 60782 205618 60866 205854
rect 61102 205618 61134 205854
rect 60514 170174 61134 205618
rect 60514 169938 60546 170174
rect 60782 169938 60866 170174
rect 61102 169938 61134 170174
rect 60514 169854 61134 169938
rect 60514 169618 60546 169854
rect 60782 169618 60866 169854
rect 61102 169618 61134 169854
rect 60514 134174 61134 169618
rect 60514 133938 60546 134174
rect 60782 133938 60866 134174
rect 61102 133938 61134 134174
rect 60514 133854 61134 133938
rect 60514 133618 60546 133854
rect 60782 133618 60866 133854
rect 61102 133618 61134 133854
rect 60514 98174 61134 133618
rect 60514 97938 60546 98174
rect 60782 97938 60866 98174
rect 61102 97938 61134 98174
rect 60514 97854 61134 97938
rect 60514 97618 60546 97854
rect 60782 97618 60866 97854
rect 61102 97618 61134 97854
rect 60514 62174 61134 97618
rect 60514 61938 60546 62174
rect 60782 61938 60866 62174
rect 61102 61938 61134 62174
rect 60514 61854 61134 61938
rect 60514 61618 60546 61854
rect 60782 61618 60866 61854
rect 61102 61618 61134 61854
rect 60514 26174 61134 61618
rect 60514 25938 60546 26174
rect 60782 25938 60866 26174
rect 61102 25938 61134 26174
rect 60514 25854 61134 25938
rect 60514 25618 60546 25854
rect 60782 25618 60866 25854
rect 61102 25618 61134 25854
rect 57838 3229 57898 11782
rect 57835 3228 57901 3229
rect 57835 3164 57836 3228
rect 57900 3164 57901 3228
rect 57835 3163 57901 3164
rect 56794 -5382 56826 -5146
rect 57062 -5382 57146 -5146
rect 57382 -5382 57414 -5146
rect 56794 -5466 57414 -5382
rect 56794 -5702 56826 -5466
rect 57062 -5702 57146 -5466
rect 57382 -5702 57414 -5466
rect 56794 -7654 57414 -5702
rect 60514 -6106 61134 25618
rect 60514 -6342 60546 -6106
rect 60782 -6342 60866 -6106
rect 61102 -6342 61134 -6106
rect 60514 -6426 61134 -6342
rect 60514 -6662 60546 -6426
rect 60782 -6662 60866 -6426
rect 61102 -6662 61134 -6426
rect 60514 -7654 61134 -6662
rect 64234 711558 64854 711590
rect 64234 711322 64266 711558
rect 64502 711322 64586 711558
rect 64822 711322 64854 711558
rect 64234 711238 64854 711322
rect 64234 711002 64266 711238
rect 64502 711002 64586 711238
rect 64822 711002 64854 711238
rect 64234 677894 64854 711002
rect 64234 677658 64266 677894
rect 64502 677658 64586 677894
rect 64822 677658 64854 677894
rect 64234 677574 64854 677658
rect 64234 677338 64266 677574
rect 64502 677338 64586 677574
rect 64822 677338 64854 677574
rect 64234 641894 64854 677338
rect 64234 641658 64266 641894
rect 64502 641658 64586 641894
rect 64822 641658 64854 641894
rect 64234 641574 64854 641658
rect 64234 641338 64266 641574
rect 64502 641338 64586 641574
rect 64822 641338 64854 641574
rect 64234 605894 64854 641338
rect 64234 605658 64266 605894
rect 64502 605658 64586 605894
rect 64822 605658 64854 605894
rect 64234 605574 64854 605658
rect 64234 605338 64266 605574
rect 64502 605338 64586 605574
rect 64822 605338 64854 605574
rect 64234 569894 64854 605338
rect 64234 569658 64266 569894
rect 64502 569658 64586 569894
rect 64822 569658 64854 569894
rect 64234 569574 64854 569658
rect 64234 569338 64266 569574
rect 64502 569338 64586 569574
rect 64822 569338 64854 569574
rect 64234 533894 64854 569338
rect 64234 533658 64266 533894
rect 64502 533658 64586 533894
rect 64822 533658 64854 533894
rect 64234 533574 64854 533658
rect 64234 533338 64266 533574
rect 64502 533338 64586 533574
rect 64822 533338 64854 533574
rect 64234 497894 64854 533338
rect 64234 497658 64266 497894
rect 64502 497658 64586 497894
rect 64822 497658 64854 497894
rect 64234 497574 64854 497658
rect 64234 497338 64266 497574
rect 64502 497338 64586 497574
rect 64822 497338 64854 497574
rect 64234 461894 64854 497338
rect 64234 461658 64266 461894
rect 64502 461658 64586 461894
rect 64822 461658 64854 461894
rect 64234 461574 64854 461658
rect 64234 461338 64266 461574
rect 64502 461338 64586 461574
rect 64822 461338 64854 461574
rect 64234 425894 64854 461338
rect 64234 425658 64266 425894
rect 64502 425658 64586 425894
rect 64822 425658 64854 425894
rect 64234 425574 64854 425658
rect 64234 425338 64266 425574
rect 64502 425338 64586 425574
rect 64822 425338 64854 425574
rect 64234 389894 64854 425338
rect 64234 389658 64266 389894
rect 64502 389658 64586 389894
rect 64822 389658 64854 389894
rect 64234 389574 64854 389658
rect 64234 389338 64266 389574
rect 64502 389338 64586 389574
rect 64822 389338 64854 389574
rect 64234 353894 64854 389338
rect 64234 353658 64266 353894
rect 64502 353658 64586 353894
rect 64822 353658 64854 353894
rect 64234 353574 64854 353658
rect 64234 353338 64266 353574
rect 64502 353338 64586 353574
rect 64822 353338 64854 353574
rect 64234 317894 64854 353338
rect 64234 317658 64266 317894
rect 64502 317658 64586 317894
rect 64822 317658 64854 317894
rect 64234 317574 64854 317658
rect 64234 317338 64266 317574
rect 64502 317338 64586 317574
rect 64822 317338 64854 317574
rect 64234 281894 64854 317338
rect 64234 281658 64266 281894
rect 64502 281658 64586 281894
rect 64822 281658 64854 281894
rect 64234 281574 64854 281658
rect 64234 281338 64266 281574
rect 64502 281338 64586 281574
rect 64822 281338 64854 281574
rect 64234 245894 64854 281338
rect 64234 245658 64266 245894
rect 64502 245658 64586 245894
rect 64822 245658 64854 245894
rect 64234 245574 64854 245658
rect 64234 245338 64266 245574
rect 64502 245338 64586 245574
rect 64822 245338 64854 245574
rect 64234 209894 64854 245338
rect 64234 209658 64266 209894
rect 64502 209658 64586 209894
rect 64822 209658 64854 209894
rect 64234 209574 64854 209658
rect 64234 209338 64266 209574
rect 64502 209338 64586 209574
rect 64822 209338 64854 209574
rect 64234 173894 64854 209338
rect 64234 173658 64266 173894
rect 64502 173658 64586 173894
rect 64822 173658 64854 173894
rect 64234 173574 64854 173658
rect 64234 173338 64266 173574
rect 64502 173338 64586 173574
rect 64822 173338 64854 173574
rect 64234 137894 64854 173338
rect 64234 137658 64266 137894
rect 64502 137658 64586 137894
rect 64822 137658 64854 137894
rect 64234 137574 64854 137658
rect 64234 137338 64266 137574
rect 64502 137338 64586 137574
rect 64822 137338 64854 137574
rect 64234 101894 64854 137338
rect 64234 101658 64266 101894
rect 64502 101658 64586 101894
rect 64822 101658 64854 101894
rect 64234 101574 64854 101658
rect 64234 101338 64266 101574
rect 64502 101338 64586 101574
rect 64822 101338 64854 101574
rect 64234 65894 64854 101338
rect 64234 65658 64266 65894
rect 64502 65658 64586 65894
rect 64822 65658 64854 65894
rect 64234 65574 64854 65658
rect 64234 65338 64266 65574
rect 64502 65338 64586 65574
rect 64822 65338 64854 65574
rect 64234 29894 64854 65338
rect 64234 29658 64266 29894
rect 64502 29658 64586 29894
rect 64822 29658 64854 29894
rect 64234 29574 64854 29658
rect 64234 29338 64266 29574
rect 64502 29338 64586 29574
rect 64822 29338 64854 29574
rect 64234 -7066 64854 29338
rect 74194 704838 74814 711590
rect 74194 704602 74226 704838
rect 74462 704602 74546 704838
rect 74782 704602 74814 704838
rect 74194 704518 74814 704602
rect 74194 704282 74226 704518
rect 74462 704282 74546 704518
rect 74782 704282 74814 704518
rect 74194 687854 74814 704282
rect 74194 687618 74226 687854
rect 74462 687618 74546 687854
rect 74782 687618 74814 687854
rect 74194 687534 74814 687618
rect 74194 687298 74226 687534
rect 74462 687298 74546 687534
rect 74782 687298 74814 687534
rect 74194 651854 74814 687298
rect 74194 651618 74226 651854
rect 74462 651618 74546 651854
rect 74782 651618 74814 651854
rect 74194 651534 74814 651618
rect 74194 651298 74226 651534
rect 74462 651298 74546 651534
rect 74782 651298 74814 651534
rect 74194 615854 74814 651298
rect 74194 615618 74226 615854
rect 74462 615618 74546 615854
rect 74782 615618 74814 615854
rect 74194 615534 74814 615618
rect 74194 615298 74226 615534
rect 74462 615298 74546 615534
rect 74782 615298 74814 615534
rect 74194 579854 74814 615298
rect 74194 579618 74226 579854
rect 74462 579618 74546 579854
rect 74782 579618 74814 579854
rect 74194 579534 74814 579618
rect 74194 579298 74226 579534
rect 74462 579298 74546 579534
rect 74782 579298 74814 579534
rect 74194 543854 74814 579298
rect 74194 543618 74226 543854
rect 74462 543618 74546 543854
rect 74782 543618 74814 543854
rect 74194 543534 74814 543618
rect 74194 543298 74226 543534
rect 74462 543298 74546 543534
rect 74782 543298 74814 543534
rect 74194 507854 74814 543298
rect 74194 507618 74226 507854
rect 74462 507618 74546 507854
rect 74782 507618 74814 507854
rect 74194 507534 74814 507618
rect 74194 507298 74226 507534
rect 74462 507298 74546 507534
rect 74782 507298 74814 507534
rect 74194 471854 74814 507298
rect 74194 471618 74226 471854
rect 74462 471618 74546 471854
rect 74782 471618 74814 471854
rect 74194 471534 74814 471618
rect 74194 471298 74226 471534
rect 74462 471298 74546 471534
rect 74782 471298 74814 471534
rect 74194 435854 74814 471298
rect 74194 435618 74226 435854
rect 74462 435618 74546 435854
rect 74782 435618 74814 435854
rect 74194 435534 74814 435618
rect 74194 435298 74226 435534
rect 74462 435298 74546 435534
rect 74782 435298 74814 435534
rect 74194 399854 74814 435298
rect 74194 399618 74226 399854
rect 74462 399618 74546 399854
rect 74782 399618 74814 399854
rect 74194 399534 74814 399618
rect 74194 399298 74226 399534
rect 74462 399298 74546 399534
rect 74782 399298 74814 399534
rect 74194 363854 74814 399298
rect 74194 363618 74226 363854
rect 74462 363618 74546 363854
rect 74782 363618 74814 363854
rect 74194 363534 74814 363618
rect 74194 363298 74226 363534
rect 74462 363298 74546 363534
rect 74782 363298 74814 363534
rect 74194 327854 74814 363298
rect 74194 327618 74226 327854
rect 74462 327618 74546 327854
rect 74782 327618 74814 327854
rect 74194 327534 74814 327618
rect 74194 327298 74226 327534
rect 74462 327298 74546 327534
rect 74782 327298 74814 327534
rect 74194 291854 74814 327298
rect 74194 291618 74226 291854
rect 74462 291618 74546 291854
rect 74782 291618 74814 291854
rect 74194 291534 74814 291618
rect 74194 291298 74226 291534
rect 74462 291298 74546 291534
rect 74782 291298 74814 291534
rect 74194 255854 74814 291298
rect 74194 255618 74226 255854
rect 74462 255618 74546 255854
rect 74782 255618 74814 255854
rect 74194 255534 74814 255618
rect 74194 255298 74226 255534
rect 74462 255298 74546 255534
rect 74782 255298 74814 255534
rect 74194 219854 74814 255298
rect 74194 219618 74226 219854
rect 74462 219618 74546 219854
rect 74782 219618 74814 219854
rect 74194 219534 74814 219618
rect 74194 219298 74226 219534
rect 74462 219298 74546 219534
rect 74782 219298 74814 219534
rect 74194 183854 74814 219298
rect 74194 183618 74226 183854
rect 74462 183618 74546 183854
rect 74782 183618 74814 183854
rect 74194 183534 74814 183618
rect 74194 183298 74226 183534
rect 74462 183298 74546 183534
rect 74782 183298 74814 183534
rect 74194 147854 74814 183298
rect 74194 147618 74226 147854
rect 74462 147618 74546 147854
rect 74782 147618 74814 147854
rect 74194 147534 74814 147618
rect 74194 147298 74226 147534
rect 74462 147298 74546 147534
rect 74782 147298 74814 147534
rect 74194 111854 74814 147298
rect 74194 111618 74226 111854
rect 74462 111618 74546 111854
rect 74782 111618 74814 111854
rect 74194 111534 74814 111618
rect 74194 111298 74226 111534
rect 74462 111298 74546 111534
rect 74782 111298 74814 111534
rect 74194 75854 74814 111298
rect 74194 75618 74226 75854
rect 74462 75618 74546 75854
rect 74782 75618 74814 75854
rect 74194 75534 74814 75618
rect 74194 75298 74226 75534
rect 74462 75298 74546 75534
rect 74782 75298 74814 75534
rect 74194 39854 74814 75298
rect 74194 39618 74226 39854
rect 74462 39618 74546 39854
rect 74782 39618 74814 39854
rect 74194 39534 74814 39618
rect 74194 39298 74226 39534
rect 74462 39298 74546 39534
rect 74782 39298 74814 39534
rect 67406 3229 67466 8382
rect 70347 5948 70413 5949
rect 70347 5884 70348 5948
rect 70412 5884 70413 5948
rect 70347 5883 70413 5884
rect 70350 3229 70410 5883
rect 74194 3854 74814 39298
rect 77914 705798 78534 711590
rect 77914 705562 77946 705798
rect 78182 705562 78266 705798
rect 78502 705562 78534 705798
rect 77914 705478 78534 705562
rect 77914 705242 77946 705478
rect 78182 705242 78266 705478
rect 78502 705242 78534 705478
rect 77914 691574 78534 705242
rect 77914 691338 77946 691574
rect 78182 691338 78266 691574
rect 78502 691338 78534 691574
rect 77914 691254 78534 691338
rect 77914 691018 77946 691254
rect 78182 691018 78266 691254
rect 78502 691018 78534 691254
rect 77914 655574 78534 691018
rect 77914 655338 77946 655574
rect 78182 655338 78266 655574
rect 78502 655338 78534 655574
rect 77914 655254 78534 655338
rect 77914 655018 77946 655254
rect 78182 655018 78266 655254
rect 78502 655018 78534 655254
rect 77914 619574 78534 655018
rect 77914 619338 77946 619574
rect 78182 619338 78266 619574
rect 78502 619338 78534 619574
rect 77914 619254 78534 619338
rect 77914 619018 77946 619254
rect 78182 619018 78266 619254
rect 78502 619018 78534 619254
rect 77914 583574 78534 619018
rect 77914 583338 77946 583574
rect 78182 583338 78266 583574
rect 78502 583338 78534 583574
rect 77914 583254 78534 583338
rect 77914 583018 77946 583254
rect 78182 583018 78266 583254
rect 78502 583018 78534 583254
rect 77914 547574 78534 583018
rect 77914 547338 77946 547574
rect 78182 547338 78266 547574
rect 78502 547338 78534 547574
rect 77914 547254 78534 547338
rect 77914 547018 77946 547254
rect 78182 547018 78266 547254
rect 78502 547018 78534 547254
rect 77914 511574 78534 547018
rect 77914 511338 77946 511574
rect 78182 511338 78266 511574
rect 78502 511338 78534 511574
rect 77914 511254 78534 511338
rect 77914 511018 77946 511254
rect 78182 511018 78266 511254
rect 78502 511018 78534 511254
rect 77914 475574 78534 511018
rect 77914 475338 77946 475574
rect 78182 475338 78266 475574
rect 78502 475338 78534 475574
rect 77914 475254 78534 475338
rect 77914 475018 77946 475254
rect 78182 475018 78266 475254
rect 78502 475018 78534 475254
rect 77914 439574 78534 475018
rect 77914 439338 77946 439574
rect 78182 439338 78266 439574
rect 78502 439338 78534 439574
rect 77914 439254 78534 439338
rect 77914 439018 77946 439254
rect 78182 439018 78266 439254
rect 78502 439018 78534 439254
rect 77914 403574 78534 439018
rect 77914 403338 77946 403574
rect 78182 403338 78266 403574
rect 78502 403338 78534 403574
rect 77914 403254 78534 403338
rect 77914 403018 77946 403254
rect 78182 403018 78266 403254
rect 78502 403018 78534 403254
rect 77914 367574 78534 403018
rect 77914 367338 77946 367574
rect 78182 367338 78266 367574
rect 78502 367338 78534 367574
rect 77914 367254 78534 367338
rect 77914 367018 77946 367254
rect 78182 367018 78266 367254
rect 78502 367018 78534 367254
rect 77914 331574 78534 367018
rect 77914 331338 77946 331574
rect 78182 331338 78266 331574
rect 78502 331338 78534 331574
rect 77914 331254 78534 331338
rect 77914 331018 77946 331254
rect 78182 331018 78266 331254
rect 78502 331018 78534 331254
rect 77914 295574 78534 331018
rect 77914 295338 77946 295574
rect 78182 295338 78266 295574
rect 78502 295338 78534 295574
rect 77914 295254 78534 295338
rect 77914 295018 77946 295254
rect 78182 295018 78266 295254
rect 78502 295018 78534 295254
rect 77914 259574 78534 295018
rect 77914 259338 77946 259574
rect 78182 259338 78266 259574
rect 78502 259338 78534 259574
rect 77914 259254 78534 259338
rect 77914 259018 77946 259254
rect 78182 259018 78266 259254
rect 78502 259018 78534 259254
rect 77914 223574 78534 259018
rect 77914 223338 77946 223574
rect 78182 223338 78266 223574
rect 78502 223338 78534 223574
rect 77914 223254 78534 223338
rect 77914 223018 77946 223254
rect 78182 223018 78266 223254
rect 78502 223018 78534 223254
rect 77914 187574 78534 223018
rect 77914 187338 77946 187574
rect 78182 187338 78266 187574
rect 78502 187338 78534 187574
rect 77914 187254 78534 187338
rect 77914 187018 77946 187254
rect 78182 187018 78266 187254
rect 78502 187018 78534 187254
rect 77914 151574 78534 187018
rect 77914 151338 77946 151574
rect 78182 151338 78266 151574
rect 78502 151338 78534 151574
rect 77914 151254 78534 151338
rect 77914 151018 77946 151254
rect 78182 151018 78266 151254
rect 78502 151018 78534 151254
rect 77914 115574 78534 151018
rect 77914 115338 77946 115574
rect 78182 115338 78266 115574
rect 78502 115338 78534 115574
rect 77914 115254 78534 115338
rect 77914 115018 77946 115254
rect 78182 115018 78266 115254
rect 78502 115018 78534 115254
rect 77914 79574 78534 115018
rect 77914 79338 77946 79574
rect 78182 79338 78266 79574
rect 78502 79338 78534 79574
rect 77914 79254 78534 79338
rect 77914 79018 77946 79254
rect 78182 79018 78266 79254
rect 78502 79018 78534 79254
rect 77914 43574 78534 79018
rect 77914 43338 77946 43574
rect 78182 43338 78266 43574
rect 78502 43338 78534 43574
rect 77914 43254 78534 43338
rect 77914 43018 77946 43254
rect 78182 43018 78266 43254
rect 78502 43018 78534 43254
rect 77339 7852 77405 7853
rect 77339 7850 77340 7852
rect 77158 7790 77340 7850
rect 77158 6085 77218 7790
rect 77339 7788 77340 7790
rect 77404 7788 77405 7852
rect 77339 7787 77405 7788
rect 77914 7574 78534 43018
rect 77914 7338 77946 7574
rect 78182 7338 78266 7574
rect 78502 7338 78534 7574
rect 77914 7254 78534 7338
rect 77914 7018 77946 7254
rect 78182 7018 78266 7254
rect 78502 7018 78534 7254
rect 77155 6084 77221 6085
rect 77155 6020 77156 6084
rect 77220 6020 77221 6084
rect 77155 6019 77221 6020
rect 74194 3618 74226 3854
rect 74462 3618 74546 3854
rect 74782 3618 74814 3854
rect 74194 3534 74814 3618
rect 74194 3298 74226 3534
rect 74462 3298 74546 3534
rect 74782 3298 74814 3534
rect 67403 3228 67469 3229
rect 67403 3164 67404 3228
rect 67468 3164 67469 3228
rect 67403 3163 67469 3164
rect 70347 3228 70413 3229
rect 70347 3164 70348 3228
rect 70412 3164 70413 3228
rect 70347 3163 70413 3164
rect 64234 -7302 64266 -7066
rect 64502 -7302 64586 -7066
rect 64822 -7302 64854 -7066
rect 64234 -7386 64854 -7302
rect 64234 -7622 64266 -7386
rect 64502 -7622 64586 -7386
rect 64822 -7622 64854 -7386
rect 64234 -7654 64854 -7622
rect 74194 -346 74814 3298
rect 74194 -582 74226 -346
rect 74462 -582 74546 -346
rect 74782 -582 74814 -346
rect 74194 -666 74814 -582
rect 74194 -902 74226 -666
rect 74462 -902 74546 -666
rect 74782 -902 74814 -666
rect 74194 -7654 74814 -902
rect 77914 -1306 78534 7018
rect 77914 -1542 77946 -1306
rect 78182 -1542 78266 -1306
rect 78502 -1542 78534 -1306
rect 77914 -1626 78534 -1542
rect 77914 -1862 77946 -1626
rect 78182 -1862 78266 -1626
rect 78502 -1862 78534 -1626
rect 77914 -7654 78534 -1862
rect 81634 706758 82254 711590
rect 81634 706522 81666 706758
rect 81902 706522 81986 706758
rect 82222 706522 82254 706758
rect 81634 706438 82254 706522
rect 81634 706202 81666 706438
rect 81902 706202 81986 706438
rect 82222 706202 82254 706438
rect 81634 695294 82254 706202
rect 81634 695058 81666 695294
rect 81902 695058 81986 695294
rect 82222 695058 82254 695294
rect 81634 694974 82254 695058
rect 81634 694738 81666 694974
rect 81902 694738 81986 694974
rect 82222 694738 82254 694974
rect 81634 659294 82254 694738
rect 81634 659058 81666 659294
rect 81902 659058 81986 659294
rect 82222 659058 82254 659294
rect 81634 658974 82254 659058
rect 81634 658738 81666 658974
rect 81902 658738 81986 658974
rect 82222 658738 82254 658974
rect 81634 623294 82254 658738
rect 81634 623058 81666 623294
rect 81902 623058 81986 623294
rect 82222 623058 82254 623294
rect 81634 622974 82254 623058
rect 81634 622738 81666 622974
rect 81902 622738 81986 622974
rect 82222 622738 82254 622974
rect 81634 587294 82254 622738
rect 81634 587058 81666 587294
rect 81902 587058 81986 587294
rect 82222 587058 82254 587294
rect 81634 586974 82254 587058
rect 81634 586738 81666 586974
rect 81902 586738 81986 586974
rect 82222 586738 82254 586974
rect 81634 551294 82254 586738
rect 81634 551058 81666 551294
rect 81902 551058 81986 551294
rect 82222 551058 82254 551294
rect 81634 550974 82254 551058
rect 81634 550738 81666 550974
rect 81902 550738 81986 550974
rect 82222 550738 82254 550974
rect 81634 515294 82254 550738
rect 81634 515058 81666 515294
rect 81902 515058 81986 515294
rect 82222 515058 82254 515294
rect 81634 514974 82254 515058
rect 81634 514738 81666 514974
rect 81902 514738 81986 514974
rect 82222 514738 82254 514974
rect 81634 479294 82254 514738
rect 81634 479058 81666 479294
rect 81902 479058 81986 479294
rect 82222 479058 82254 479294
rect 81634 478974 82254 479058
rect 81634 478738 81666 478974
rect 81902 478738 81986 478974
rect 82222 478738 82254 478974
rect 81634 443294 82254 478738
rect 81634 443058 81666 443294
rect 81902 443058 81986 443294
rect 82222 443058 82254 443294
rect 81634 442974 82254 443058
rect 81634 442738 81666 442974
rect 81902 442738 81986 442974
rect 82222 442738 82254 442974
rect 81634 407294 82254 442738
rect 81634 407058 81666 407294
rect 81902 407058 81986 407294
rect 82222 407058 82254 407294
rect 81634 406974 82254 407058
rect 81634 406738 81666 406974
rect 81902 406738 81986 406974
rect 82222 406738 82254 406974
rect 81634 371294 82254 406738
rect 81634 371058 81666 371294
rect 81902 371058 81986 371294
rect 82222 371058 82254 371294
rect 81634 370974 82254 371058
rect 81634 370738 81666 370974
rect 81902 370738 81986 370974
rect 82222 370738 82254 370974
rect 81634 335294 82254 370738
rect 81634 335058 81666 335294
rect 81902 335058 81986 335294
rect 82222 335058 82254 335294
rect 81634 334974 82254 335058
rect 81634 334738 81666 334974
rect 81902 334738 81986 334974
rect 82222 334738 82254 334974
rect 81634 299294 82254 334738
rect 81634 299058 81666 299294
rect 81902 299058 81986 299294
rect 82222 299058 82254 299294
rect 81634 298974 82254 299058
rect 81634 298738 81666 298974
rect 81902 298738 81986 298974
rect 82222 298738 82254 298974
rect 81634 263294 82254 298738
rect 81634 263058 81666 263294
rect 81902 263058 81986 263294
rect 82222 263058 82254 263294
rect 81634 262974 82254 263058
rect 81634 262738 81666 262974
rect 81902 262738 81986 262974
rect 82222 262738 82254 262974
rect 81634 227294 82254 262738
rect 81634 227058 81666 227294
rect 81902 227058 81986 227294
rect 82222 227058 82254 227294
rect 81634 226974 82254 227058
rect 81634 226738 81666 226974
rect 81902 226738 81986 226974
rect 82222 226738 82254 226974
rect 81634 191294 82254 226738
rect 81634 191058 81666 191294
rect 81902 191058 81986 191294
rect 82222 191058 82254 191294
rect 81634 190974 82254 191058
rect 81634 190738 81666 190974
rect 81902 190738 81986 190974
rect 82222 190738 82254 190974
rect 81634 155294 82254 190738
rect 85354 707718 85974 711590
rect 85354 707482 85386 707718
rect 85622 707482 85706 707718
rect 85942 707482 85974 707718
rect 85354 707398 85974 707482
rect 85354 707162 85386 707398
rect 85622 707162 85706 707398
rect 85942 707162 85974 707398
rect 85354 699014 85974 707162
rect 85354 698778 85386 699014
rect 85622 698778 85706 699014
rect 85942 698778 85974 699014
rect 85354 698694 85974 698778
rect 85354 698458 85386 698694
rect 85622 698458 85706 698694
rect 85942 698458 85974 698694
rect 85354 663014 85974 698458
rect 85354 662778 85386 663014
rect 85622 662778 85706 663014
rect 85942 662778 85974 663014
rect 85354 662694 85974 662778
rect 85354 662458 85386 662694
rect 85622 662458 85706 662694
rect 85942 662458 85974 662694
rect 85354 627014 85974 662458
rect 85354 626778 85386 627014
rect 85622 626778 85706 627014
rect 85942 626778 85974 627014
rect 85354 626694 85974 626778
rect 85354 626458 85386 626694
rect 85622 626458 85706 626694
rect 85942 626458 85974 626694
rect 85354 591014 85974 626458
rect 85354 590778 85386 591014
rect 85622 590778 85706 591014
rect 85942 590778 85974 591014
rect 85354 590694 85974 590778
rect 85354 590458 85386 590694
rect 85622 590458 85706 590694
rect 85942 590458 85974 590694
rect 85354 555014 85974 590458
rect 85354 554778 85386 555014
rect 85622 554778 85706 555014
rect 85942 554778 85974 555014
rect 85354 554694 85974 554778
rect 85354 554458 85386 554694
rect 85622 554458 85706 554694
rect 85942 554458 85974 554694
rect 85354 519014 85974 554458
rect 85354 518778 85386 519014
rect 85622 518778 85706 519014
rect 85942 518778 85974 519014
rect 85354 518694 85974 518778
rect 85354 518458 85386 518694
rect 85622 518458 85706 518694
rect 85942 518458 85974 518694
rect 85354 483014 85974 518458
rect 85354 482778 85386 483014
rect 85622 482778 85706 483014
rect 85942 482778 85974 483014
rect 85354 482694 85974 482778
rect 85354 482458 85386 482694
rect 85622 482458 85706 482694
rect 85942 482458 85974 482694
rect 85354 447014 85974 482458
rect 85354 446778 85386 447014
rect 85622 446778 85706 447014
rect 85942 446778 85974 447014
rect 85354 446694 85974 446778
rect 85354 446458 85386 446694
rect 85622 446458 85706 446694
rect 85942 446458 85974 446694
rect 85354 411014 85974 446458
rect 85354 410778 85386 411014
rect 85622 410778 85706 411014
rect 85942 410778 85974 411014
rect 85354 410694 85974 410778
rect 85354 410458 85386 410694
rect 85622 410458 85706 410694
rect 85942 410458 85974 410694
rect 85354 375014 85974 410458
rect 85354 374778 85386 375014
rect 85622 374778 85706 375014
rect 85942 374778 85974 375014
rect 85354 374694 85974 374778
rect 85354 374458 85386 374694
rect 85622 374458 85706 374694
rect 85942 374458 85974 374694
rect 85354 339014 85974 374458
rect 85354 338778 85386 339014
rect 85622 338778 85706 339014
rect 85942 338778 85974 339014
rect 85354 338694 85974 338778
rect 85354 338458 85386 338694
rect 85622 338458 85706 338694
rect 85942 338458 85974 338694
rect 85354 303014 85974 338458
rect 85354 302778 85386 303014
rect 85622 302778 85706 303014
rect 85942 302778 85974 303014
rect 85354 302694 85974 302778
rect 85354 302458 85386 302694
rect 85622 302458 85706 302694
rect 85942 302458 85974 302694
rect 85354 267014 85974 302458
rect 85354 266778 85386 267014
rect 85622 266778 85706 267014
rect 85942 266778 85974 267014
rect 85354 266694 85974 266778
rect 85354 266458 85386 266694
rect 85622 266458 85706 266694
rect 85942 266458 85974 266694
rect 85354 231014 85974 266458
rect 85354 230778 85386 231014
rect 85622 230778 85706 231014
rect 85942 230778 85974 231014
rect 85354 230694 85974 230778
rect 85354 230458 85386 230694
rect 85622 230458 85706 230694
rect 85942 230458 85974 230694
rect 85354 195014 85974 230458
rect 85354 194778 85386 195014
rect 85622 194778 85706 195014
rect 85942 194778 85974 195014
rect 85354 194694 85974 194778
rect 85354 194458 85386 194694
rect 85622 194458 85706 194694
rect 85942 194458 85974 194694
rect 84208 183854 84528 183886
rect 84208 183618 84250 183854
rect 84486 183618 84528 183854
rect 84208 183534 84528 183618
rect 84208 183298 84250 183534
rect 84486 183298 84528 183534
rect 84208 183266 84528 183298
rect 81634 155058 81666 155294
rect 81902 155058 81986 155294
rect 82222 155058 82254 155294
rect 81634 154974 82254 155058
rect 81634 154738 81666 154974
rect 81902 154738 81986 154974
rect 82222 154738 82254 154974
rect 81634 119294 82254 154738
rect 85354 159014 85974 194458
rect 85354 158778 85386 159014
rect 85622 158778 85706 159014
rect 85942 158778 85974 159014
rect 85354 158694 85974 158778
rect 85354 158458 85386 158694
rect 85622 158458 85706 158694
rect 85942 158458 85974 158694
rect 84208 147854 84528 147886
rect 84208 147618 84250 147854
rect 84486 147618 84528 147854
rect 84208 147534 84528 147618
rect 84208 147298 84250 147534
rect 84486 147298 84528 147534
rect 84208 147266 84528 147298
rect 81634 119058 81666 119294
rect 81902 119058 81986 119294
rect 82222 119058 82254 119294
rect 81634 118974 82254 119058
rect 81634 118738 81666 118974
rect 81902 118738 81986 118974
rect 82222 118738 82254 118974
rect 81634 83294 82254 118738
rect 85354 123014 85974 158458
rect 85354 122778 85386 123014
rect 85622 122778 85706 123014
rect 85942 122778 85974 123014
rect 85354 122694 85974 122778
rect 85354 122458 85386 122694
rect 85622 122458 85706 122694
rect 85942 122458 85974 122694
rect 84208 111854 84528 111886
rect 84208 111618 84250 111854
rect 84486 111618 84528 111854
rect 84208 111534 84528 111618
rect 84208 111298 84250 111534
rect 84486 111298 84528 111534
rect 84208 111266 84528 111298
rect 81634 83058 81666 83294
rect 81902 83058 81986 83294
rect 82222 83058 82254 83294
rect 81634 82974 82254 83058
rect 81634 82738 81666 82974
rect 81902 82738 81986 82974
rect 82222 82738 82254 82974
rect 81634 47294 82254 82738
rect 81634 47058 81666 47294
rect 81902 47058 81986 47294
rect 82222 47058 82254 47294
rect 81634 46974 82254 47058
rect 81634 46738 81666 46974
rect 81902 46738 81986 46974
rect 82222 46738 82254 46974
rect 81634 11294 82254 46738
rect 81634 11058 81666 11294
rect 81902 11058 81986 11294
rect 82222 11058 82254 11294
rect 81634 10974 82254 11058
rect 81634 10738 81666 10974
rect 81902 10738 81986 10974
rect 82222 10738 82254 10974
rect 81634 -2266 82254 10738
rect 81634 -2502 81666 -2266
rect 81902 -2502 81986 -2266
rect 82222 -2502 82254 -2266
rect 81634 -2586 82254 -2502
rect 81634 -2822 81666 -2586
rect 81902 -2822 81986 -2586
rect 82222 -2822 82254 -2586
rect 81634 -7654 82254 -2822
rect 85354 87014 85974 122458
rect 85354 86778 85386 87014
rect 85622 86778 85706 87014
rect 85942 86778 85974 87014
rect 85354 86694 85974 86778
rect 85354 86458 85386 86694
rect 85622 86458 85706 86694
rect 85942 86458 85974 86694
rect 85354 51014 85974 86458
rect 85354 50778 85386 51014
rect 85622 50778 85706 51014
rect 85942 50778 85974 51014
rect 85354 50694 85974 50778
rect 85354 50458 85386 50694
rect 85622 50458 85706 50694
rect 85942 50458 85974 50694
rect 85354 15014 85974 50458
rect 85354 14778 85386 15014
rect 85622 14778 85706 15014
rect 85942 14778 85974 15014
rect 85354 14694 85974 14778
rect 85354 14458 85386 14694
rect 85622 14458 85706 14694
rect 85942 14458 85974 14694
rect 85354 -3226 85974 14458
rect 85354 -3462 85386 -3226
rect 85622 -3462 85706 -3226
rect 85942 -3462 85974 -3226
rect 85354 -3546 85974 -3462
rect 85354 -3782 85386 -3546
rect 85622 -3782 85706 -3546
rect 85942 -3782 85974 -3546
rect 85354 -7654 85974 -3782
rect 89074 708678 89694 711590
rect 89074 708442 89106 708678
rect 89342 708442 89426 708678
rect 89662 708442 89694 708678
rect 89074 708358 89694 708442
rect 89074 708122 89106 708358
rect 89342 708122 89426 708358
rect 89662 708122 89694 708358
rect 89074 666734 89694 708122
rect 89074 666498 89106 666734
rect 89342 666498 89426 666734
rect 89662 666498 89694 666734
rect 89074 666414 89694 666498
rect 89074 666178 89106 666414
rect 89342 666178 89426 666414
rect 89662 666178 89694 666414
rect 89074 630734 89694 666178
rect 89074 630498 89106 630734
rect 89342 630498 89426 630734
rect 89662 630498 89694 630734
rect 89074 630414 89694 630498
rect 89074 630178 89106 630414
rect 89342 630178 89426 630414
rect 89662 630178 89694 630414
rect 89074 594734 89694 630178
rect 89074 594498 89106 594734
rect 89342 594498 89426 594734
rect 89662 594498 89694 594734
rect 89074 594414 89694 594498
rect 89074 594178 89106 594414
rect 89342 594178 89426 594414
rect 89662 594178 89694 594414
rect 89074 558734 89694 594178
rect 89074 558498 89106 558734
rect 89342 558498 89426 558734
rect 89662 558498 89694 558734
rect 89074 558414 89694 558498
rect 89074 558178 89106 558414
rect 89342 558178 89426 558414
rect 89662 558178 89694 558414
rect 89074 522734 89694 558178
rect 89074 522498 89106 522734
rect 89342 522498 89426 522734
rect 89662 522498 89694 522734
rect 89074 522414 89694 522498
rect 89074 522178 89106 522414
rect 89342 522178 89426 522414
rect 89662 522178 89694 522414
rect 89074 486734 89694 522178
rect 89074 486498 89106 486734
rect 89342 486498 89426 486734
rect 89662 486498 89694 486734
rect 89074 486414 89694 486498
rect 89074 486178 89106 486414
rect 89342 486178 89426 486414
rect 89662 486178 89694 486414
rect 89074 450734 89694 486178
rect 89074 450498 89106 450734
rect 89342 450498 89426 450734
rect 89662 450498 89694 450734
rect 89074 450414 89694 450498
rect 89074 450178 89106 450414
rect 89342 450178 89426 450414
rect 89662 450178 89694 450414
rect 89074 414734 89694 450178
rect 89074 414498 89106 414734
rect 89342 414498 89426 414734
rect 89662 414498 89694 414734
rect 89074 414414 89694 414498
rect 89074 414178 89106 414414
rect 89342 414178 89426 414414
rect 89662 414178 89694 414414
rect 89074 378734 89694 414178
rect 89074 378498 89106 378734
rect 89342 378498 89426 378734
rect 89662 378498 89694 378734
rect 89074 378414 89694 378498
rect 89074 378178 89106 378414
rect 89342 378178 89426 378414
rect 89662 378178 89694 378414
rect 89074 342734 89694 378178
rect 89074 342498 89106 342734
rect 89342 342498 89426 342734
rect 89662 342498 89694 342734
rect 89074 342414 89694 342498
rect 89074 342178 89106 342414
rect 89342 342178 89426 342414
rect 89662 342178 89694 342414
rect 89074 306734 89694 342178
rect 89074 306498 89106 306734
rect 89342 306498 89426 306734
rect 89662 306498 89694 306734
rect 89074 306414 89694 306498
rect 89074 306178 89106 306414
rect 89342 306178 89426 306414
rect 89662 306178 89694 306414
rect 89074 270734 89694 306178
rect 89074 270498 89106 270734
rect 89342 270498 89426 270734
rect 89662 270498 89694 270734
rect 89074 270414 89694 270498
rect 89074 270178 89106 270414
rect 89342 270178 89426 270414
rect 89662 270178 89694 270414
rect 89074 234734 89694 270178
rect 89074 234498 89106 234734
rect 89342 234498 89426 234734
rect 89662 234498 89694 234734
rect 89074 234414 89694 234498
rect 89074 234178 89106 234414
rect 89342 234178 89426 234414
rect 89662 234178 89694 234414
rect 89074 198734 89694 234178
rect 89074 198498 89106 198734
rect 89342 198498 89426 198734
rect 89662 198498 89694 198734
rect 89074 198414 89694 198498
rect 89074 198178 89106 198414
rect 89342 198178 89426 198414
rect 89662 198178 89694 198414
rect 89074 162734 89694 198178
rect 89074 162498 89106 162734
rect 89342 162498 89426 162734
rect 89662 162498 89694 162734
rect 89074 162414 89694 162498
rect 89074 162178 89106 162414
rect 89342 162178 89426 162414
rect 89662 162178 89694 162414
rect 89074 126734 89694 162178
rect 89074 126498 89106 126734
rect 89342 126498 89426 126734
rect 89662 126498 89694 126734
rect 89074 126414 89694 126498
rect 89074 126178 89106 126414
rect 89342 126178 89426 126414
rect 89662 126178 89694 126414
rect 89074 90734 89694 126178
rect 89074 90498 89106 90734
rect 89342 90498 89426 90734
rect 89662 90498 89694 90734
rect 89074 90414 89694 90498
rect 89074 90178 89106 90414
rect 89342 90178 89426 90414
rect 89662 90178 89694 90414
rect 89074 54734 89694 90178
rect 92794 709638 93414 711590
rect 92794 709402 92826 709638
rect 93062 709402 93146 709638
rect 93382 709402 93414 709638
rect 92794 709318 93414 709402
rect 92794 709082 92826 709318
rect 93062 709082 93146 709318
rect 93382 709082 93414 709318
rect 92794 670454 93414 709082
rect 92794 670218 92826 670454
rect 93062 670218 93146 670454
rect 93382 670218 93414 670454
rect 92794 670134 93414 670218
rect 92794 669898 92826 670134
rect 93062 669898 93146 670134
rect 93382 669898 93414 670134
rect 92794 634454 93414 669898
rect 92794 634218 92826 634454
rect 93062 634218 93146 634454
rect 93382 634218 93414 634454
rect 92794 634134 93414 634218
rect 92794 633898 92826 634134
rect 93062 633898 93146 634134
rect 93382 633898 93414 634134
rect 92794 598454 93414 633898
rect 92794 598218 92826 598454
rect 93062 598218 93146 598454
rect 93382 598218 93414 598454
rect 92794 598134 93414 598218
rect 92794 597898 92826 598134
rect 93062 597898 93146 598134
rect 93382 597898 93414 598134
rect 92794 562454 93414 597898
rect 92794 562218 92826 562454
rect 93062 562218 93146 562454
rect 93382 562218 93414 562454
rect 92794 562134 93414 562218
rect 92794 561898 92826 562134
rect 93062 561898 93146 562134
rect 93382 561898 93414 562134
rect 92794 526454 93414 561898
rect 92794 526218 92826 526454
rect 93062 526218 93146 526454
rect 93382 526218 93414 526454
rect 92794 526134 93414 526218
rect 92794 525898 92826 526134
rect 93062 525898 93146 526134
rect 93382 525898 93414 526134
rect 92794 490454 93414 525898
rect 92794 490218 92826 490454
rect 93062 490218 93146 490454
rect 93382 490218 93414 490454
rect 92794 490134 93414 490218
rect 92794 489898 92826 490134
rect 93062 489898 93146 490134
rect 93382 489898 93414 490134
rect 92794 454454 93414 489898
rect 92794 454218 92826 454454
rect 93062 454218 93146 454454
rect 93382 454218 93414 454454
rect 92794 454134 93414 454218
rect 92794 453898 92826 454134
rect 93062 453898 93146 454134
rect 93382 453898 93414 454134
rect 92794 418454 93414 453898
rect 92794 418218 92826 418454
rect 93062 418218 93146 418454
rect 93382 418218 93414 418454
rect 92794 418134 93414 418218
rect 92794 417898 92826 418134
rect 93062 417898 93146 418134
rect 93382 417898 93414 418134
rect 92794 382454 93414 417898
rect 92794 382218 92826 382454
rect 93062 382218 93146 382454
rect 93382 382218 93414 382454
rect 92794 382134 93414 382218
rect 92794 381898 92826 382134
rect 93062 381898 93146 382134
rect 93382 381898 93414 382134
rect 92794 346454 93414 381898
rect 92794 346218 92826 346454
rect 93062 346218 93146 346454
rect 93382 346218 93414 346454
rect 92794 346134 93414 346218
rect 92794 345898 92826 346134
rect 93062 345898 93146 346134
rect 93382 345898 93414 346134
rect 92794 310454 93414 345898
rect 92794 310218 92826 310454
rect 93062 310218 93146 310454
rect 93382 310218 93414 310454
rect 92794 310134 93414 310218
rect 92794 309898 92826 310134
rect 93062 309898 93146 310134
rect 93382 309898 93414 310134
rect 92794 274454 93414 309898
rect 92794 274218 92826 274454
rect 93062 274218 93146 274454
rect 93382 274218 93414 274454
rect 92794 274134 93414 274218
rect 92794 273898 92826 274134
rect 93062 273898 93146 274134
rect 93382 273898 93414 274134
rect 92794 238454 93414 273898
rect 92794 238218 92826 238454
rect 93062 238218 93146 238454
rect 93382 238218 93414 238454
rect 92794 238134 93414 238218
rect 92794 237898 92826 238134
rect 93062 237898 93146 238134
rect 93382 237898 93414 238134
rect 92794 202454 93414 237898
rect 92794 202218 92826 202454
rect 93062 202218 93146 202454
rect 93382 202218 93414 202454
rect 92794 202134 93414 202218
rect 92794 201898 92826 202134
rect 93062 201898 93146 202134
rect 93382 201898 93414 202134
rect 92794 166454 93414 201898
rect 92794 166218 92826 166454
rect 93062 166218 93146 166454
rect 93382 166218 93414 166454
rect 92794 166134 93414 166218
rect 92794 165898 92826 166134
rect 93062 165898 93146 166134
rect 93382 165898 93414 166134
rect 92794 130454 93414 165898
rect 92794 130218 92826 130454
rect 93062 130218 93146 130454
rect 93382 130218 93414 130454
rect 92794 130134 93414 130218
rect 92794 129898 92826 130134
rect 93062 129898 93146 130134
rect 93382 129898 93414 130134
rect 92794 94454 93414 129898
rect 92794 94218 92826 94454
rect 93062 94218 93146 94454
rect 93382 94218 93414 94454
rect 92794 94134 93414 94218
rect 92794 93898 92826 94134
rect 93062 93898 93146 94134
rect 93382 93898 93414 94134
rect 91139 77348 91205 77349
rect 91139 77284 91140 77348
rect 91204 77284 91205 77348
rect 91139 77283 91205 77284
rect 89074 54498 89106 54734
rect 89342 54498 89426 54734
rect 89662 54498 89694 54734
rect 89074 54414 89694 54498
rect 89074 54178 89106 54414
rect 89342 54178 89426 54414
rect 89662 54178 89694 54414
rect 89074 18734 89694 54178
rect 89074 18498 89106 18734
rect 89342 18498 89426 18734
rect 89662 18498 89694 18734
rect 89074 18414 89694 18498
rect 89074 18178 89106 18414
rect 89342 18178 89426 18414
rect 89662 18178 89694 18414
rect 89074 -4186 89694 18178
rect 91142 4538 91202 77283
rect 92794 58454 93414 93898
rect 96514 710598 97134 711590
rect 96514 710362 96546 710598
rect 96782 710362 96866 710598
rect 97102 710362 97134 710598
rect 96514 710278 97134 710362
rect 96514 710042 96546 710278
rect 96782 710042 96866 710278
rect 97102 710042 97134 710278
rect 96514 674174 97134 710042
rect 96514 673938 96546 674174
rect 96782 673938 96866 674174
rect 97102 673938 97134 674174
rect 96514 673854 97134 673938
rect 96514 673618 96546 673854
rect 96782 673618 96866 673854
rect 97102 673618 97134 673854
rect 96514 638174 97134 673618
rect 96514 637938 96546 638174
rect 96782 637938 96866 638174
rect 97102 637938 97134 638174
rect 96514 637854 97134 637938
rect 96514 637618 96546 637854
rect 96782 637618 96866 637854
rect 97102 637618 97134 637854
rect 96514 602174 97134 637618
rect 96514 601938 96546 602174
rect 96782 601938 96866 602174
rect 97102 601938 97134 602174
rect 96514 601854 97134 601938
rect 96514 601618 96546 601854
rect 96782 601618 96866 601854
rect 97102 601618 97134 601854
rect 96514 566174 97134 601618
rect 96514 565938 96546 566174
rect 96782 565938 96866 566174
rect 97102 565938 97134 566174
rect 96514 565854 97134 565938
rect 96514 565618 96546 565854
rect 96782 565618 96866 565854
rect 97102 565618 97134 565854
rect 96514 530174 97134 565618
rect 96514 529938 96546 530174
rect 96782 529938 96866 530174
rect 97102 529938 97134 530174
rect 96514 529854 97134 529938
rect 96514 529618 96546 529854
rect 96782 529618 96866 529854
rect 97102 529618 97134 529854
rect 96514 494174 97134 529618
rect 96514 493938 96546 494174
rect 96782 493938 96866 494174
rect 97102 493938 97134 494174
rect 96514 493854 97134 493938
rect 96514 493618 96546 493854
rect 96782 493618 96866 493854
rect 97102 493618 97134 493854
rect 96514 458174 97134 493618
rect 96514 457938 96546 458174
rect 96782 457938 96866 458174
rect 97102 457938 97134 458174
rect 96514 457854 97134 457938
rect 96514 457618 96546 457854
rect 96782 457618 96866 457854
rect 97102 457618 97134 457854
rect 96514 422174 97134 457618
rect 96514 421938 96546 422174
rect 96782 421938 96866 422174
rect 97102 421938 97134 422174
rect 96514 421854 97134 421938
rect 96514 421618 96546 421854
rect 96782 421618 96866 421854
rect 97102 421618 97134 421854
rect 96514 386174 97134 421618
rect 96514 385938 96546 386174
rect 96782 385938 96866 386174
rect 97102 385938 97134 386174
rect 96514 385854 97134 385938
rect 96514 385618 96546 385854
rect 96782 385618 96866 385854
rect 97102 385618 97134 385854
rect 96514 350174 97134 385618
rect 96514 349938 96546 350174
rect 96782 349938 96866 350174
rect 97102 349938 97134 350174
rect 96514 349854 97134 349938
rect 96514 349618 96546 349854
rect 96782 349618 96866 349854
rect 97102 349618 97134 349854
rect 96514 314174 97134 349618
rect 96514 313938 96546 314174
rect 96782 313938 96866 314174
rect 97102 313938 97134 314174
rect 96514 313854 97134 313938
rect 96514 313618 96546 313854
rect 96782 313618 96866 313854
rect 97102 313618 97134 313854
rect 96514 278174 97134 313618
rect 96514 277938 96546 278174
rect 96782 277938 96866 278174
rect 97102 277938 97134 278174
rect 96514 277854 97134 277938
rect 96514 277618 96546 277854
rect 96782 277618 96866 277854
rect 97102 277618 97134 277854
rect 96514 242174 97134 277618
rect 96514 241938 96546 242174
rect 96782 241938 96866 242174
rect 97102 241938 97134 242174
rect 96514 241854 97134 241938
rect 96514 241618 96546 241854
rect 96782 241618 96866 241854
rect 97102 241618 97134 241854
rect 96514 206174 97134 241618
rect 96514 205938 96546 206174
rect 96782 205938 96866 206174
rect 97102 205938 97134 206174
rect 96514 205854 97134 205938
rect 96514 205618 96546 205854
rect 96782 205618 96866 205854
rect 97102 205618 97134 205854
rect 96514 170174 97134 205618
rect 100234 711558 100854 711590
rect 100234 711322 100266 711558
rect 100502 711322 100586 711558
rect 100822 711322 100854 711558
rect 100234 711238 100854 711322
rect 100234 711002 100266 711238
rect 100502 711002 100586 711238
rect 100822 711002 100854 711238
rect 100234 677894 100854 711002
rect 100234 677658 100266 677894
rect 100502 677658 100586 677894
rect 100822 677658 100854 677894
rect 100234 677574 100854 677658
rect 100234 677338 100266 677574
rect 100502 677338 100586 677574
rect 100822 677338 100854 677574
rect 100234 641894 100854 677338
rect 100234 641658 100266 641894
rect 100502 641658 100586 641894
rect 100822 641658 100854 641894
rect 100234 641574 100854 641658
rect 100234 641338 100266 641574
rect 100502 641338 100586 641574
rect 100822 641338 100854 641574
rect 100234 605894 100854 641338
rect 100234 605658 100266 605894
rect 100502 605658 100586 605894
rect 100822 605658 100854 605894
rect 100234 605574 100854 605658
rect 100234 605338 100266 605574
rect 100502 605338 100586 605574
rect 100822 605338 100854 605574
rect 100234 569894 100854 605338
rect 100234 569658 100266 569894
rect 100502 569658 100586 569894
rect 100822 569658 100854 569894
rect 100234 569574 100854 569658
rect 100234 569338 100266 569574
rect 100502 569338 100586 569574
rect 100822 569338 100854 569574
rect 100234 533894 100854 569338
rect 100234 533658 100266 533894
rect 100502 533658 100586 533894
rect 100822 533658 100854 533894
rect 100234 533574 100854 533658
rect 100234 533338 100266 533574
rect 100502 533338 100586 533574
rect 100822 533338 100854 533574
rect 100234 497894 100854 533338
rect 100234 497658 100266 497894
rect 100502 497658 100586 497894
rect 100822 497658 100854 497894
rect 100234 497574 100854 497658
rect 100234 497338 100266 497574
rect 100502 497338 100586 497574
rect 100822 497338 100854 497574
rect 100234 461894 100854 497338
rect 100234 461658 100266 461894
rect 100502 461658 100586 461894
rect 100822 461658 100854 461894
rect 100234 461574 100854 461658
rect 100234 461338 100266 461574
rect 100502 461338 100586 461574
rect 100822 461338 100854 461574
rect 100234 425894 100854 461338
rect 100234 425658 100266 425894
rect 100502 425658 100586 425894
rect 100822 425658 100854 425894
rect 100234 425574 100854 425658
rect 100234 425338 100266 425574
rect 100502 425338 100586 425574
rect 100822 425338 100854 425574
rect 100234 389894 100854 425338
rect 100234 389658 100266 389894
rect 100502 389658 100586 389894
rect 100822 389658 100854 389894
rect 100234 389574 100854 389658
rect 100234 389338 100266 389574
rect 100502 389338 100586 389574
rect 100822 389338 100854 389574
rect 100234 353894 100854 389338
rect 100234 353658 100266 353894
rect 100502 353658 100586 353894
rect 100822 353658 100854 353894
rect 100234 353574 100854 353658
rect 100234 353338 100266 353574
rect 100502 353338 100586 353574
rect 100822 353338 100854 353574
rect 100234 317894 100854 353338
rect 100234 317658 100266 317894
rect 100502 317658 100586 317894
rect 100822 317658 100854 317894
rect 100234 317574 100854 317658
rect 100234 317338 100266 317574
rect 100502 317338 100586 317574
rect 100822 317338 100854 317574
rect 100234 281894 100854 317338
rect 100234 281658 100266 281894
rect 100502 281658 100586 281894
rect 100822 281658 100854 281894
rect 100234 281574 100854 281658
rect 100234 281338 100266 281574
rect 100502 281338 100586 281574
rect 100822 281338 100854 281574
rect 100234 245894 100854 281338
rect 100234 245658 100266 245894
rect 100502 245658 100586 245894
rect 100822 245658 100854 245894
rect 100234 245574 100854 245658
rect 100234 245338 100266 245574
rect 100502 245338 100586 245574
rect 100822 245338 100854 245574
rect 100234 209894 100854 245338
rect 100234 209658 100266 209894
rect 100502 209658 100586 209894
rect 100822 209658 100854 209894
rect 100234 209574 100854 209658
rect 100234 209338 100266 209574
rect 100502 209338 100586 209574
rect 100822 209338 100854 209574
rect 100234 188457 100854 209338
rect 110194 704838 110814 711590
rect 110194 704602 110226 704838
rect 110462 704602 110546 704838
rect 110782 704602 110814 704838
rect 110194 704518 110814 704602
rect 110194 704282 110226 704518
rect 110462 704282 110546 704518
rect 110782 704282 110814 704518
rect 110194 687854 110814 704282
rect 110194 687618 110226 687854
rect 110462 687618 110546 687854
rect 110782 687618 110814 687854
rect 110194 687534 110814 687618
rect 110194 687298 110226 687534
rect 110462 687298 110546 687534
rect 110782 687298 110814 687534
rect 110194 651854 110814 687298
rect 110194 651618 110226 651854
rect 110462 651618 110546 651854
rect 110782 651618 110814 651854
rect 110194 651534 110814 651618
rect 110194 651298 110226 651534
rect 110462 651298 110546 651534
rect 110782 651298 110814 651534
rect 110194 615854 110814 651298
rect 110194 615618 110226 615854
rect 110462 615618 110546 615854
rect 110782 615618 110814 615854
rect 110194 615534 110814 615618
rect 110194 615298 110226 615534
rect 110462 615298 110546 615534
rect 110782 615298 110814 615534
rect 110194 579854 110814 615298
rect 110194 579618 110226 579854
rect 110462 579618 110546 579854
rect 110782 579618 110814 579854
rect 110194 579534 110814 579618
rect 110194 579298 110226 579534
rect 110462 579298 110546 579534
rect 110782 579298 110814 579534
rect 110194 543854 110814 579298
rect 110194 543618 110226 543854
rect 110462 543618 110546 543854
rect 110782 543618 110814 543854
rect 110194 543534 110814 543618
rect 110194 543298 110226 543534
rect 110462 543298 110546 543534
rect 110782 543298 110814 543534
rect 110194 507854 110814 543298
rect 110194 507618 110226 507854
rect 110462 507618 110546 507854
rect 110782 507618 110814 507854
rect 110194 507534 110814 507618
rect 110194 507298 110226 507534
rect 110462 507298 110546 507534
rect 110782 507298 110814 507534
rect 110194 471854 110814 507298
rect 110194 471618 110226 471854
rect 110462 471618 110546 471854
rect 110782 471618 110814 471854
rect 110194 471534 110814 471618
rect 110194 471298 110226 471534
rect 110462 471298 110546 471534
rect 110782 471298 110814 471534
rect 110194 435854 110814 471298
rect 110194 435618 110226 435854
rect 110462 435618 110546 435854
rect 110782 435618 110814 435854
rect 110194 435534 110814 435618
rect 110194 435298 110226 435534
rect 110462 435298 110546 435534
rect 110782 435298 110814 435534
rect 110194 399854 110814 435298
rect 110194 399618 110226 399854
rect 110462 399618 110546 399854
rect 110782 399618 110814 399854
rect 110194 399534 110814 399618
rect 110194 399298 110226 399534
rect 110462 399298 110546 399534
rect 110782 399298 110814 399534
rect 110194 363854 110814 399298
rect 110194 363618 110226 363854
rect 110462 363618 110546 363854
rect 110782 363618 110814 363854
rect 110194 363534 110814 363618
rect 110194 363298 110226 363534
rect 110462 363298 110546 363534
rect 110782 363298 110814 363534
rect 110194 327854 110814 363298
rect 110194 327618 110226 327854
rect 110462 327618 110546 327854
rect 110782 327618 110814 327854
rect 110194 327534 110814 327618
rect 110194 327298 110226 327534
rect 110462 327298 110546 327534
rect 110782 327298 110814 327534
rect 110194 291854 110814 327298
rect 110194 291618 110226 291854
rect 110462 291618 110546 291854
rect 110782 291618 110814 291854
rect 110194 291534 110814 291618
rect 110194 291298 110226 291534
rect 110462 291298 110546 291534
rect 110782 291298 110814 291534
rect 110194 255854 110814 291298
rect 110194 255618 110226 255854
rect 110462 255618 110546 255854
rect 110782 255618 110814 255854
rect 110194 255534 110814 255618
rect 110194 255298 110226 255534
rect 110462 255298 110546 255534
rect 110782 255298 110814 255534
rect 110194 219854 110814 255298
rect 110194 219618 110226 219854
rect 110462 219618 110546 219854
rect 110782 219618 110814 219854
rect 110194 219534 110814 219618
rect 110194 219298 110226 219534
rect 110462 219298 110546 219534
rect 110782 219298 110814 219534
rect 110194 188457 110814 219298
rect 113914 705798 114534 711590
rect 113914 705562 113946 705798
rect 114182 705562 114266 705798
rect 114502 705562 114534 705798
rect 113914 705478 114534 705562
rect 113914 705242 113946 705478
rect 114182 705242 114266 705478
rect 114502 705242 114534 705478
rect 113914 691574 114534 705242
rect 113914 691338 113946 691574
rect 114182 691338 114266 691574
rect 114502 691338 114534 691574
rect 113914 691254 114534 691338
rect 113914 691018 113946 691254
rect 114182 691018 114266 691254
rect 114502 691018 114534 691254
rect 113914 655574 114534 691018
rect 113914 655338 113946 655574
rect 114182 655338 114266 655574
rect 114502 655338 114534 655574
rect 113914 655254 114534 655338
rect 113914 655018 113946 655254
rect 114182 655018 114266 655254
rect 114502 655018 114534 655254
rect 113914 619574 114534 655018
rect 113914 619338 113946 619574
rect 114182 619338 114266 619574
rect 114502 619338 114534 619574
rect 113914 619254 114534 619338
rect 113914 619018 113946 619254
rect 114182 619018 114266 619254
rect 114502 619018 114534 619254
rect 113914 583574 114534 619018
rect 113914 583338 113946 583574
rect 114182 583338 114266 583574
rect 114502 583338 114534 583574
rect 113914 583254 114534 583338
rect 113914 583018 113946 583254
rect 114182 583018 114266 583254
rect 114502 583018 114534 583254
rect 113914 547574 114534 583018
rect 113914 547338 113946 547574
rect 114182 547338 114266 547574
rect 114502 547338 114534 547574
rect 113914 547254 114534 547338
rect 113914 547018 113946 547254
rect 114182 547018 114266 547254
rect 114502 547018 114534 547254
rect 113914 511574 114534 547018
rect 113914 511338 113946 511574
rect 114182 511338 114266 511574
rect 114502 511338 114534 511574
rect 113914 511254 114534 511338
rect 113914 511018 113946 511254
rect 114182 511018 114266 511254
rect 114502 511018 114534 511254
rect 113914 475574 114534 511018
rect 113914 475338 113946 475574
rect 114182 475338 114266 475574
rect 114502 475338 114534 475574
rect 113914 475254 114534 475338
rect 113914 475018 113946 475254
rect 114182 475018 114266 475254
rect 114502 475018 114534 475254
rect 113914 439574 114534 475018
rect 113914 439338 113946 439574
rect 114182 439338 114266 439574
rect 114502 439338 114534 439574
rect 113914 439254 114534 439338
rect 113914 439018 113946 439254
rect 114182 439018 114266 439254
rect 114502 439018 114534 439254
rect 113914 403574 114534 439018
rect 113914 403338 113946 403574
rect 114182 403338 114266 403574
rect 114502 403338 114534 403574
rect 113914 403254 114534 403338
rect 113914 403018 113946 403254
rect 114182 403018 114266 403254
rect 114502 403018 114534 403254
rect 113914 367574 114534 403018
rect 113914 367338 113946 367574
rect 114182 367338 114266 367574
rect 114502 367338 114534 367574
rect 113914 367254 114534 367338
rect 113914 367018 113946 367254
rect 114182 367018 114266 367254
rect 114502 367018 114534 367254
rect 113914 331574 114534 367018
rect 113914 331338 113946 331574
rect 114182 331338 114266 331574
rect 114502 331338 114534 331574
rect 113914 331254 114534 331338
rect 113914 331018 113946 331254
rect 114182 331018 114266 331254
rect 114502 331018 114534 331254
rect 113914 295574 114534 331018
rect 113914 295338 113946 295574
rect 114182 295338 114266 295574
rect 114502 295338 114534 295574
rect 113914 295254 114534 295338
rect 113914 295018 113946 295254
rect 114182 295018 114266 295254
rect 114502 295018 114534 295254
rect 113914 259574 114534 295018
rect 113914 259338 113946 259574
rect 114182 259338 114266 259574
rect 114502 259338 114534 259574
rect 113914 259254 114534 259338
rect 113914 259018 113946 259254
rect 114182 259018 114266 259254
rect 114502 259018 114534 259254
rect 113914 223574 114534 259018
rect 113914 223338 113946 223574
rect 114182 223338 114266 223574
rect 114502 223338 114534 223574
rect 113914 223254 114534 223338
rect 113914 223018 113946 223254
rect 114182 223018 114266 223254
rect 114502 223018 114534 223254
rect 113914 188457 114534 223018
rect 117634 706758 118254 711590
rect 117634 706522 117666 706758
rect 117902 706522 117986 706758
rect 118222 706522 118254 706758
rect 117634 706438 118254 706522
rect 117634 706202 117666 706438
rect 117902 706202 117986 706438
rect 118222 706202 118254 706438
rect 117634 695294 118254 706202
rect 117634 695058 117666 695294
rect 117902 695058 117986 695294
rect 118222 695058 118254 695294
rect 117634 694974 118254 695058
rect 117634 694738 117666 694974
rect 117902 694738 117986 694974
rect 118222 694738 118254 694974
rect 117634 659294 118254 694738
rect 117634 659058 117666 659294
rect 117902 659058 117986 659294
rect 118222 659058 118254 659294
rect 117634 658974 118254 659058
rect 117634 658738 117666 658974
rect 117902 658738 117986 658974
rect 118222 658738 118254 658974
rect 117634 623294 118254 658738
rect 117634 623058 117666 623294
rect 117902 623058 117986 623294
rect 118222 623058 118254 623294
rect 117634 622974 118254 623058
rect 117634 622738 117666 622974
rect 117902 622738 117986 622974
rect 118222 622738 118254 622974
rect 117634 587294 118254 622738
rect 117634 587058 117666 587294
rect 117902 587058 117986 587294
rect 118222 587058 118254 587294
rect 117634 586974 118254 587058
rect 117634 586738 117666 586974
rect 117902 586738 117986 586974
rect 118222 586738 118254 586974
rect 117634 551294 118254 586738
rect 117634 551058 117666 551294
rect 117902 551058 117986 551294
rect 118222 551058 118254 551294
rect 117634 550974 118254 551058
rect 117634 550738 117666 550974
rect 117902 550738 117986 550974
rect 118222 550738 118254 550974
rect 117634 515294 118254 550738
rect 117634 515058 117666 515294
rect 117902 515058 117986 515294
rect 118222 515058 118254 515294
rect 117634 514974 118254 515058
rect 117634 514738 117666 514974
rect 117902 514738 117986 514974
rect 118222 514738 118254 514974
rect 117634 479294 118254 514738
rect 117634 479058 117666 479294
rect 117902 479058 117986 479294
rect 118222 479058 118254 479294
rect 117634 478974 118254 479058
rect 117634 478738 117666 478974
rect 117902 478738 117986 478974
rect 118222 478738 118254 478974
rect 117634 443294 118254 478738
rect 117634 443058 117666 443294
rect 117902 443058 117986 443294
rect 118222 443058 118254 443294
rect 117634 442974 118254 443058
rect 117634 442738 117666 442974
rect 117902 442738 117986 442974
rect 118222 442738 118254 442974
rect 117634 407294 118254 442738
rect 117634 407058 117666 407294
rect 117902 407058 117986 407294
rect 118222 407058 118254 407294
rect 117634 406974 118254 407058
rect 117634 406738 117666 406974
rect 117902 406738 117986 406974
rect 118222 406738 118254 406974
rect 117634 371294 118254 406738
rect 117634 371058 117666 371294
rect 117902 371058 117986 371294
rect 118222 371058 118254 371294
rect 117634 370974 118254 371058
rect 117634 370738 117666 370974
rect 117902 370738 117986 370974
rect 118222 370738 118254 370974
rect 117634 335294 118254 370738
rect 117634 335058 117666 335294
rect 117902 335058 117986 335294
rect 118222 335058 118254 335294
rect 117634 334974 118254 335058
rect 117634 334738 117666 334974
rect 117902 334738 117986 334974
rect 118222 334738 118254 334974
rect 117634 299294 118254 334738
rect 117634 299058 117666 299294
rect 117902 299058 117986 299294
rect 118222 299058 118254 299294
rect 117634 298974 118254 299058
rect 117634 298738 117666 298974
rect 117902 298738 117986 298974
rect 118222 298738 118254 298974
rect 117634 263294 118254 298738
rect 117634 263058 117666 263294
rect 117902 263058 117986 263294
rect 118222 263058 118254 263294
rect 117634 262974 118254 263058
rect 117634 262738 117666 262974
rect 117902 262738 117986 262974
rect 118222 262738 118254 262974
rect 117634 227294 118254 262738
rect 117634 227058 117666 227294
rect 117902 227058 117986 227294
rect 118222 227058 118254 227294
rect 117634 226974 118254 227058
rect 117634 226738 117666 226974
rect 117902 226738 117986 226974
rect 118222 226738 118254 226974
rect 117634 191294 118254 226738
rect 117634 191058 117666 191294
rect 117902 191058 117986 191294
rect 118222 191058 118254 191294
rect 117634 190974 118254 191058
rect 117634 190738 117666 190974
rect 117902 190738 117986 190974
rect 118222 190738 118254 190974
rect 117634 188457 118254 190738
rect 121354 707718 121974 711590
rect 121354 707482 121386 707718
rect 121622 707482 121706 707718
rect 121942 707482 121974 707718
rect 121354 707398 121974 707482
rect 121354 707162 121386 707398
rect 121622 707162 121706 707398
rect 121942 707162 121974 707398
rect 121354 699014 121974 707162
rect 121354 698778 121386 699014
rect 121622 698778 121706 699014
rect 121942 698778 121974 699014
rect 121354 698694 121974 698778
rect 121354 698458 121386 698694
rect 121622 698458 121706 698694
rect 121942 698458 121974 698694
rect 121354 663014 121974 698458
rect 121354 662778 121386 663014
rect 121622 662778 121706 663014
rect 121942 662778 121974 663014
rect 121354 662694 121974 662778
rect 121354 662458 121386 662694
rect 121622 662458 121706 662694
rect 121942 662458 121974 662694
rect 121354 627014 121974 662458
rect 121354 626778 121386 627014
rect 121622 626778 121706 627014
rect 121942 626778 121974 627014
rect 121354 626694 121974 626778
rect 121354 626458 121386 626694
rect 121622 626458 121706 626694
rect 121942 626458 121974 626694
rect 121354 591014 121974 626458
rect 121354 590778 121386 591014
rect 121622 590778 121706 591014
rect 121942 590778 121974 591014
rect 121354 590694 121974 590778
rect 121354 590458 121386 590694
rect 121622 590458 121706 590694
rect 121942 590458 121974 590694
rect 121354 555014 121974 590458
rect 121354 554778 121386 555014
rect 121622 554778 121706 555014
rect 121942 554778 121974 555014
rect 121354 554694 121974 554778
rect 121354 554458 121386 554694
rect 121622 554458 121706 554694
rect 121942 554458 121974 554694
rect 121354 519014 121974 554458
rect 121354 518778 121386 519014
rect 121622 518778 121706 519014
rect 121942 518778 121974 519014
rect 121354 518694 121974 518778
rect 121354 518458 121386 518694
rect 121622 518458 121706 518694
rect 121942 518458 121974 518694
rect 121354 483014 121974 518458
rect 121354 482778 121386 483014
rect 121622 482778 121706 483014
rect 121942 482778 121974 483014
rect 121354 482694 121974 482778
rect 121354 482458 121386 482694
rect 121622 482458 121706 482694
rect 121942 482458 121974 482694
rect 121354 447014 121974 482458
rect 121354 446778 121386 447014
rect 121622 446778 121706 447014
rect 121942 446778 121974 447014
rect 121354 446694 121974 446778
rect 121354 446458 121386 446694
rect 121622 446458 121706 446694
rect 121942 446458 121974 446694
rect 121354 411014 121974 446458
rect 121354 410778 121386 411014
rect 121622 410778 121706 411014
rect 121942 410778 121974 411014
rect 121354 410694 121974 410778
rect 121354 410458 121386 410694
rect 121622 410458 121706 410694
rect 121942 410458 121974 410694
rect 121354 375014 121974 410458
rect 121354 374778 121386 375014
rect 121622 374778 121706 375014
rect 121942 374778 121974 375014
rect 121354 374694 121974 374778
rect 121354 374458 121386 374694
rect 121622 374458 121706 374694
rect 121942 374458 121974 374694
rect 121354 339014 121974 374458
rect 121354 338778 121386 339014
rect 121622 338778 121706 339014
rect 121942 338778 121974 339014
rect 121354 338694 121974 338778
rect 121354 338458 121386 338694
rect 121622 338458 121706 338694
rect 121942 338458 121974 338694
rect 121354 303014 121974 338458
rect 121354 302778 121386 303014
rect 121622 302778 121706 303014
rect 121942 302778 121974 303014
rect 121354 302694 121974 302778
rect 121354 302458 121386 302694
rect 121622 302458 121706 302694
rect 121942 302458 121974 302694
rect 121354 267014 121974 302458
rect 121354 266778 121386 267014
rect 121622 266778 121706 267014
rect 121942 266778 121974 267014
rect 121354 266694 121974 266778
rect 121354 266458 121386 266694
rect 121622 266458 121706 266694
rect 121942 266458 121974 266694
rect 121354 231014 121974 266458
rect 121354 230778 121386 231014
rect 121622 230778 121706 231014
rect 121942 230778 121974 231014
rect 121354 230694 121974 230778
rect 121354 230458 121386 230694
rect 121622 230458 121706 230694
rect 121942 230458 121974 230694
rect 121354 195014 121974 230458
rect 121354 194778 121386 195014
rect 121622 194778 121706 195014
rect 121942 194778 121974 195014
rect 121354 194694 121974 194778
rect 121354 194458 121386 194694
rect 121622 194458 121706 194694
rect 121942 194458 121974 194694
rect 121354 188457 121974 194458
rect 125074 708678 125694 711590
rect 125074 708442 125106 708678
rect 125342 708442 125426 708678
rect 125662 708442 125694 708678
rect 125074 708358 125694 708442
rect 125074 708122 125106 708358
rect 125342 708122 125426 708358
rect 125662 708122 125694 708358
rect 125074 666734 125694 708122
rect 125074 666498 125106 666734
rect 125342 666498 125426 666734
rect 125662 666498 125694 666734
rect 125074 666414 125694 666498
rect 125074 666178 125106 666414
rect 125342 666178 125426 666414
rect 125662 666178 125694 666414
rect 125074 630734 125694 666178
rect 125074 630498 125106 630734
rect 125342 630498 125426 630734
rect 125662 630498 125694 630734
rect 125074 630414 125694 630498
rect 125074 630178 125106 630414
rect 125342 630178 125426 630414
rect 125662 630178 125694 630414
rect 125074 594734 125694 630178
rect 125074 594498 125106 594734
rect 125342 594498 125426 594734
rect 125662 594498 125694 594734
rect 125074 594414 125694 594498
rect 125074 594178 125106 594414
rect 125342 594178 125426 594414
rect 125662 594178 125694 594414
rect 125074 558734 125694 594178
rect 125074 558498 125106 558734
rect 125342 558498 125426 558734
rect 125662 558498 125694 558734
rect 125074 558414 125694 558498
rect 125074 558178 125106 558414
rect 125342 558178 125426 558414
rect 125662 558178 125694 558414
rect 125074 522734 125694 558178
rect 125074 522498 125106 522734
rect 125342 522498 125426 522734
rect 125662 522498 125694 522734
rect 125074 522414 125694 522498
rect 125074 522178 125106 522414
rect 125342 522178 125426 522414
rect 125662 522178 125694 522414
rect 125074 486734 125694 522178
rect 125074 486498 125106 486734
rect 125342 486498 125426 486734
rect 125662 486498 125694 486734
rect 125074 486414 125694 486498
rect 125074 486178 125106 486414
rect 125342 486178 125426 486414
rect 125662 486178 125694 486414
rect 125074 450734 125694 486178
rect 125074 450498 125106 450734
rect 125342 450498 125426 450734
rect 125662 450498 125694 450734
rect 125074 450414 125694 450498
rect 125074 450178 125106 450414
rect 125342 450178 125426 450414
rect 125662 450178 125694 450414
rect 125074 414734 125694 450178
rect 125074 414498 125106 414734
rect 125342 414498 125426 414734
rect 125662 414498 125694 414734
rect 125074 414414 125694 414498
rect 125074 414178 125106 414414
rect 125342 414178 125426 414414
rect 125662 414178 125694 414414
rect 125074 378734 125694 414178
rect 125074 378498 125106 378734
rect 125342 378498 125426 378734
rect 125662 378498 125694 378734
rect 125074 378414 125694 378498
rect 125074 378178 125106 378414
rect 125342 378178 125426 378414
rect 125662 378178 125694 378414
rect 125074 342734 125694 378178
rect 125074 342498 125106 342734
rect 125342 342498 125426 342734
rect 125662 342498 125694 342734
rect 125074 342414 125694 342498
rect 125074 342178 125106 342414
rect 125342 342178 125426 342414
rect 125662 342178 125694 342414
rect 125074 306734 125694 342178
rect 125074 306498 125106 306734
rect 125342 306498 125426 306734
rect 125662 306498 125694 306734
rect 125074 306414 125694 306498
rect 125074 306178 125106 306414
rect 125342 306178 125426 306414
rect 125662 306178 125694 306414
rect 125074 270734 125694 306178
rect 125074 270498 125106 270734
rect 125342 270498 125426 270734
rect 125662 270498 125694 270734
rect 125074 270414 125694 270498
rect 125074 270178 125106 270414
rect 125342 270178 125426 270414
rect 125662 270178 125694 270414
rect 125074 234734 125694 270178
rect 125074 234498 125106 234734
rect 125342 234498 125426 234734
rect 125662 234498 125694 234734
rect 125074 234414 125694 234498
rect 125074 234178 125106 234414
rect 125342 234178 125426 234414
rect 125662 234178 125694 234414
rect 125074 198734 125694 234178
rect 125074 198498 125106 198734
rect 125342 198498 125426 198734
rect 125662 198498 125694 198734
rect 125074 198414 125694 198498
rect 125074 198178 125106 198414
rect 125342 198178 125426 198414
rect 125662 198178 125694 198414
rect 125074 188457 125694 198178
rect 128794 709638 129414 711590
rect 128794 709402 128826 709638
rect 129062 709402 129146 709638
rect 129382 709402 129414 709638
rect 128794 709318 129414 709402
rect 128794 709082 128826 709318
rect 129062 709082 129146 709318
rect 129382 709082 129414 709318
rect 128794 670454 129414 709082
rect 128794 670218 128826 670454
rect 129062 670218 129146 670454
rect 129382 670218 129414 670454
rect 128794 670134 129414 670218
rect 128794 669898 128826 670134
rect 129062 669898 129146 670134
rect 129382 669898 129414 670134
rect 128794 634454 129414 669898
rect 128794 634218 128826 634454
rect 129062 634218 129146 634454
rect 129382 634218 129414 634454
rect 128794 634134 129414 634218
rect 128794 633898 128826 634134
rect 129062 633898 129146 634134
rect 129382 633898 129414 634134
rect 128794 598454 129414 633898
rect 128794 598218 128826 598454
rect 129062 598218 129146 598454
rect 129382 598218 129414 598454
rect 128794 598134 129414 598218
rect 128794 597898 128826 598134
rect 129062 597898 129146 598134
rect 129382 597898 129414 598134
rect 128794 562454 129414 597898
rect 128794 562218 128826 562454
rect 129062 562218 129146 562454
rect 129382 562218 129414 562454
rect 128794 562134 129414 562218
rect 128794 561898 128826 562134
rect 129062 561898 129146 562134
rect 129382 561898 129414 562134
rect 128794 526454 129414 561898
rect 128794 526218 128826 526454
rect 129062 526218 129146 526454
rect 129382 526218 129414 526454
rect 128794 526134 129414 526218
rect 128794 525898 128826 526134
rect 129062 525898 129146 526134
rect 129382 525898 129414 526134
rect 128794 490454 129414 525898
rect 128794 490218 128826 490454
rect 129062 490218 129146 490454
rect 129382 490218 129414 490454
rect 128794 490134 129414 490218
rect 128794 489898 128826 490134
rect 129062 489898 129146 490134
rect 129382 489898 129414 490134
rect 128794 454454 129414 489898
rect 128794 454218 128826 454454
rect 129062 454218 129146 454454
rect 129382 454218 129414 454454
rect 128794 454134 129414 454218
rect 128794 453898 128826 454134
rect 129062 453898 129146 454134
rect 129382 453898 129414 454134
rect 128794 418454 129414 453898
rect 128794 418218 128826 418454
rect 129062 418218 129146 418454
rect 129382 418218 129414 418454
rect 128794 418134 129414 418218
rect 128794 417898 128826 418134
rect 129062 417898 129146 418134
rect 129382 417898 129414 418134
rect 128794 382454 129414 417898
rect 128794 382218 128826 382454
rect 129062 382218 129146 382454
rect 129382 382218 129414 382454
rect 128794 382134 129414 382218
rect 128794 381898 128826 382134
rect 129062 381898 129146 382134
rect 129382 381898 129414 382134
rect 128794 346454 129414 381898
rect 128794 346218 128826 346454
rect 129062 346218 129146 346454
rect 129382 346218 129414 346454
rect 128794 346134 129414 346218
rect 128794 345898 128826 346134
rect 129062 345898 129146 346134
rect 129382 345898 129414 346134
rect 128794 310454 129414 345898
rect 128794 310218 128826 310454
rect 129062 310218 129146 310454
rect 129382 310218 129414 310454
rect 128794 310134 129414 310218
rect 128794 309898 128826 310134
rect 129062 309898 129146 310134
rect 129382 309898 129414 310134
rect 128794 274454 129414 309898
rect 128794 274218 128826 274454
rect 129062 274218 129146 274454
rect 129382 274218 129414 274454
rect 128794 274134 129414 274218
rect 128794 273898 128826 274134
rect 129062 273898 129146 274134
rect 129382 273898 129414 274134
rect 128794 238454 129414 273898
rect 128794 238218 128826 238454
rect 129062 238218 129146 238454
rect 129382 238218 129414 238454
rect 128794 238134 129414 238218
rect 128794 237898 128826 238134
rect 129062 237898 129146 238134
rect 129382 237898 129414 238134
rect 128794 202454 129414 237898
rect 128794 202218 128826 202454
rect 129062 202218 129146 202454
rect 129382 202218 129414 202454
rect 128794 202134 129414 202218
rect 128794 201898 128826 202134
rect 129062 201898 129146 202134
rect 129382 201898 129414 202134
rect 128794 188457 129414 201898
rect 132514 710598 133134 711590
rect 132514 710362 132546 710598
rect 132782 710362 132866 710598
rect 133102 710362 133134 710598
rect 132514 710278 133134 710362
rect 132514 710042 132546 710278
rect 132782 710042 132866 710278
rect 133102 710042 133134 710278
rect 132514 674174 133134 710042
rect 132514 673938 132546 674174
rect 132782 673938 132866 674174
rect 133102 673938 133134 674174
rect 132514 673854 133134 673938
rect 132514 673618 132546 673854
rect 132782 673618 132866 673854
rect 133102 673618 133134 673854
rect 132514 638174 133134 673618
rect 132514 637938 132546 638174
rect 132782 637938 132866 638174
rect 133102 637938 133134 638174
rect 132514 637854 133134 637938
rect 132514 637618 132546 637854
rect 132782 637618 132866 637854
rect 133102 637618 133134 637854
rect 132514 602174 133134 637618
rect 132514 601938 132546 602174
rect 132782 601938 132866 602174
rect 133102 601938 133134 602174
rect 132514 601854 133134 601938
rect 132514 601618 132546 601854
rect 132782 601618 132866 601854
rect 133102 601618 133134 601854
rect 132514 566174 133134 601618
rect 132514 565938 132546 566174
rect 132782 565938 132866 566174
rect 133102 565938 133134 566174
rect 132514 565854 133134 565938
rect 132514 565618 132546 565854
rect 132782 565618 132866 565854
rect 133102 565618 133134 565854
rect 132514 530174 133134 565618
rect 132514 529938 132546 530174
rect 132782 529938 132866 530174
rect 133102 529938 133134 530174
rect 132514 529854 133134 529938
rect 132514 529618 132546 529854
rect 132782 529618 132866 529854
rect 133102 529618 133134 529854
rect 132514 494174 133134 529618
rect 132514 493938 132546 494174
rect 132782 493938 132866 494174
rect 133102 493938 133134 494174
rect 132514 493854 133134 493938
rect 132514 493618 132546 493854
rect 132782 493618 132866 493854
rect 133102 493618 133134 493854
rect 132514 458174 133134 493618
rect 132514 457938 132546 458174
rect 132782 457938 132866 458174
rect 133102 457938 133134 458174
rect 132514 457854 133134 457938
rect 132514 457618 132546 457854
rect 132782 457618 132866 457854
rect 133102 457618 133134 457854
rect 132514 422174 133134 457618
rect 132514 421938 132546 422174
rect 132782 421938 132866 422174
rect 133102 421938 133134 422174
rect 132514 421854 133134 421938
rect 132514 421618 132546 421854
rect 132782 421618 132866 421854
rect 133102 421618 133134 421854
rect 132514 386174 133134 421618
rect 132514 385938 132546 386174
rect 132782 385938 132866 386174
rect 133102 385938 133134 386174
rect 132514 385854 133134 385938
rect 132514 385618 132546 385854
rect 132782 385618 132866 385854
rect 133102 385618 133134 385854
rect 132514 350174 133134 385618
rect 132514 349938 132546 350174
rect 132782 349938 132866 350174
rect 133102 349938 133134 350174
rect 132514 349854 133134 349938
rect 132514 349618 132546 349854
rect 132782 349618 132866 349854
rect 133102 349618 133134 349854
rect 132514 314174 133134 349618
rect 132514 313938 132546 314174
rect 132782 313938 132866 314174
rect 133102 313938 133134 314174
rect 132514 313854 133134 313938
rect 132514 313618 132546 313854
rect 132782 313618 132866 313854
rect 133102 313618 133134 313854
rect 132514 278174 133134 313618
rect 132514 277938 132546 278174
rect 132782 277938 132866 278174
rect 133102 277938 133134 278174
rect 132514 277854 133134 277938
rect 132514 277618 132546 277854
rect 132782 277618 132866 277854
rect 133102 277618 133134 277854
rect 132514 242174 133134 277618
rect 132514 241938 132546 242174
rect 132782 241938 132866 242174
rect 133102 241938 133134 242174
rect 132514 241854 133134 241938
rect 132514 241618 132546 241854
rect 132782 241618 132866 241854
rect 133102 241618 133134 241854
rect 132514 206174 133134 241618
rect 132514 205938 132546 206174
rect 132782 205938 132866 206174
rect 133102 205938 133134 206174
rect 132514 205854 133134 205938
rect 132514 205618 132546 205854
rect 132782 205618 132866 205854
rect 133102 205618 133134 205854
rect 132514 188457 133134 205618
rect 136234 711558 136854 711590
rect 136234 711322 136266 711558
rect 136502 711322 136586 711558
rect 136822 711322 136854 711558
rect 136234 711238 136854 711322
rect 136234 711002 136266 711238
rect 136502 711002 136586 711238
rect 136822 711002 136854 711238
rect 136234 677894 136854 711002
rect 136234 677658 136266 677894
rect 136502 677658 136586 677894
rect 136822 677658 136854 677894
rect 136234 677574 136854 677658
rect 136234 677338 136266 677574
rect 136502 677338 136586 677574
rect 136822 677338 136854 677574
rect 136234 641894 136854 677338
rect 136234 641658 136266 641894
rect 136502 641658 136586 641894
rect 136822 641658 136854 641894
rect 136234 641574 136854 641658
rect 136234 641338 136266 641574
rect 136502 641338 136586 641574
rect 136822 641338 136854 641574
rect 136234 605894 136854 641338
rect 136234 605658 136266 605894
rect 136502 605658 136586 605894
rect 136822 605658 136854 605894
rect 136234 605574 136854 605658
rect 136234 605338 136266 605574
rect 136502 605338 136586 605574
rect 136822 605338 136854 605574
rect 136234 569894 136854 605338
rect 136234 569658 136266 569894
rect 136502 569658 136586 569894
rect 136822 569658 136854 569894
rect 136234 569574 136854 569658
rect 136234 569338 136266 569574
rect 136502 569338 136586 569574
rect 136822 569338 136854 569574
rect 136234 533894 136854 569338
rect 136234 533658 136266 533894
rect 136502 533658 136586 533894
rect 136822 533658 136854 533894
rect 136234 533574 136854 533658
rect 136234 533338 136266 533574
rect 136502 533338 136586 533574
rect 136822 533338 136854 533574
rect 136234 497894 136854 533338
rect 136234 497658 136266 497894
rect 136502 497658 136586 497894
rect 136822 497658 136854 497894
rect 136234 497574 136854 497658
rect 136234 497338 136266 497574
rect 136502 497338 136586 497574
rect 136822 497338 136854 497574
rect 136234 461894 136854 497338
rect 136234 461658 136266 461894
rect 136502 461658 136586 461894
rect 136822 461658 136854 461894
rect 136234 461574 136854 461658
rect 136234 461338 136266 461574
rect 136502 461338 136586 461574
rect 136822 461338 136854 461574
rect 136234 425894 136854 461338
rect 136234 425658 136266 425894
rect 136502 425658 136586 425894
rect 136822 425658 136854 425894
rect 136234 425574 136854 425658
rect 136234 425338 136266 425574
rect 136502 425338 136586 425574
rect 136822 425338 136854 425574
rect 136234 389894 136854 425338
rect 136234 389658 136266 389894
rect 136502 389658 136586 389894
rect 136822 389658 136854 389894
rect 136234 389574 136854 389658
rect 136234 389338 136266 389574
rect 136502 389338 136586 389574
rect 136822 389338 136854 389574
rect 136234 353894 136854 389338
rect 136234 353658 136266 353894
rect 136502 353658 136586 353894
rect 136822 353658 136854 353894
rect 136234 353574 136854 353658
rect 136234 353338 136266 353574
rect 136502 353338 136586 353574
rect 136822 353338 136854 353574
rect 136234 317894 136854 353338
rect 136234 317658 136266 317894
rect 136502 317658 136586 317894
rect 136822 317658 136854 317894
rect 136234 317574 136854 317658
rect 136234 317338 136266 317574
rect 136502 317338 136586 317574
rect 136822 317338 136854 317574
rect 136234 281894 136854 317338
rect 136234 281658 136266 281894
rect 136502 281658 136586 281894
rect 136822 281658 136854 281894
rect 136234 281574 136854 281658
rect 136234 281338 136266 281574
rect 136502 281338 136586 281574
rect 136822 281338 136854 281574
rect 136234 245894 136854 281338
rect 136234 245658 136266 245894
rect 136502 245658 136586 245894
rect 136822 245658 136854 245894
rect 136234 245574 136854 245658
rect 136234 245338 136266 245574
rect 136502 245338 136586 245574
rect 136822 245338 136854 245574
rect 136234 209894 136854 245338
rect 136234 209658 136266 209894
rect 136502 209658 136586 209894
rect 136822 209658 136854 209894
rect 136234 209574 136854 209658
rect 136234 209338 136266 209574
rect 136502 209338 136586 209574
rect 136822 209338 136854 209574
rect 136234 188457 136854 209338
rect 146194 704838 146814 711590
rect 146194 704602 146226 704838
rect 146462 704602 146546 704838
rect 146782 704602 146814 704838
rect 146194 704518 146814 704602
rect 146194 704282 146226 704518
rect 146462 704282 146546 704518
rect 146782 704282 146814 704518
rect 146194 687854 146814 704282
rect 146194 687618 146226 687854
rect 146462 687618 146546 687854
rect 146782 687618 146814 687854
rect 146194 687534 146814 687618
rect 146194 687298 146226 687534
rect 146462 687298 146546 687534
rect 146782 687298 146814 687534
rect 146194 651854 146814 687298
rect 146194 651618 146226 651854
rect 146462 651618 146546 651854
rect 146782 651618 146814 651854
rect 146194 651534 146814 651618
rect 146194 651298 146226 651534
rect 146462 651298 146546 651534
rect 146782 651298 146814 651534
rect 146194 615854 146814 651298
rect 146194 615618 146226 615854
rect 146462 615618 146546 615854
rect 146782 615618 146814 615854
rect 146194 615534 146814 615618
rect 146194 615298 146226 615534
rect 146462 615298 146546 615534
rect 146782 615298 146814 615534
rect 146194 579854 146814 615298
rect 146194 579618 146226 579854
rect 146462 579618 146546 579854
rect 146782 579618 146814 579854
rect 146194 579534 146814 579618
rect 146194 579298 146226 579534
rect 146462 579298 146546 579534
rect 146782 579298 146814 579534
rect 146194 543854 146814 579298
rect 146194 543618 146226 543854
rect 146462 543618 146546 543854
rect 146782 543618 146814 543854
rect 146194 543534 146814 543618
rect 146194 543298 146226 543534
rect 146462 543298 146546 543534
rect 146782 543298 146814 543534
rect 146194 507854 146814 543298
rect 146194 507618 146226 507854
rect 146462 507618 146546 507854
rect 146782 507618 146814 507854
rect 146194 507534 146814 507618
rect 146194 507298 146226 507534
rect 146462 507298 146546 507534
rect 146782 507298 146814 507534
rect 146194 471854 146814 507298
rect 146194 471618 146226 471854
rect 146462 471618 146546 471854
rect 146782 471618 146814 471854
rect 146194 471534 146814 471618
rect 146194 471298 146226 471534
rect 146462 471298 146546 471534
rect 146782 471298 146814 471534
rect 146194 435854 146814 471298
rect 146194 435618 146226 435854
rect 146462 435618 146546 435854
rect 146782 435618 146814 435854
rect 146194 435534 146814 435618
rect 146194 435298 146226 435534
rect 146462 435298 146546 435534
rect 146782 435298 146814 435534
rect 146194 399854 146814 435298
rect 146194 399618 146226 399854
rect 146462 399618 146546 399854
rect 146782 399618 146814 399854
rect 146194 399534 146814 399618
rect 146194 399298 146226 399534
rect 146462 399298 146546 399534
rect 146782 399298 146814 399534
rect 146194 363854 146814 399298
rect 146194 363618 146226 363854
rect 146462 363618 146546 363854
rect 146782 363618 146814 363854
rect 146194 363534 146814 363618
rect 146194 363298 146226 363534
rect 146462 363298 146546 363534
rect 146782 363298 146814 363534
rect 146194 327854 146814 363298
rect 146194 327618 146226 327854
rect 146462 327618 146546 327854
rect 146782 327618 146814 327854
rect 146194 327534 146814 327618
rect 146194 327298 146226 327534
rect 146462 327298 146546 327534
rect 146782 327298 146814 327534
rect 146194 291854 146814 327298
rect 146194 291618 146226 291854
rect 146462 291618 146546 291854
rect 146782 291618 146814 291854
rect 146194 291534 146814 291618
rect 146194 291298 146226 291534
rect 146462 291298 146546 291534
rect 146782 291298 146814 291534
rect 146194 255854 146814 291298
rect 146194 255618 146226 255854
rect 146462 255618 146546 255854
rect 146782 255618 146814 255854
rect 146194 255534 146814 255618
rect 146194 255298 146226 255534
rect 146462 255298 146546 255534
rect 146782 255298 146814 255534
rect 146194 219854 146814 255298
rect 146194 219618 146226 219854
rect 146462 219618 146546 219854
rect 146782 219618 146814 219854
rect 146194 219534 146814 219618
rect 146194 219298 146226 219534
rect 146462 219298 146546 219534
rect 146782 219298 146814 219534
rect 146194 188457 146814 219298
rect 149914 705798 150534 711590
rect 149914 705562 149946 705798
rect 150182 705562 150266 705798
rect 150502 705562 150534 705798
rect 149914 705478 150534 705562
rect 149914 705242 149946 705478
rect 150182 705242 150266 705478
rect 150502 705242 150534 705478
rect 149914 691574 150534 705242
rect 149914 691338 149946 691574
rect 150182 691338 150266 691574
rect 150502 691338 150534 691574
rect 149914 691254 150534 691338
rect 149914 691018 149946 691254
rect 150182 691018 150266 691254
rect 150502 691018 150534 691254
rect 149914 655574 150534 691018
rect 149914 655338 149946 655574
rect 150182 655338 150266 655574
rect 150502 655338 150534 655574
rect 149914 655254 150534 655338
rect 149914 655018 149946 655254
rect 150182 655018 150266 655254
rect 150502 655018 150534 655254
rect 149914 619574 150534 655018
rect 149914 619338 149946 619574
rect 150182 619338 150266 619574
rect 150502 619338 150534 619574
rect 149914 619254 150534 619338
rect 149914 619018 149946 619254
rect 150182 619018 150266 619254
rect 150502 619018 150534 619254
rect 149914 583574 150534 619018
rect 149914 583338 149946 583574
rect 150182 583338 150266 583574
rect 150502 583338 150534 583574
rect 149914 583254 150534 583338
rect 149914 583018 149946 583254
rect 150182 583018 150266 583254
rect 150502 583018 150534 583254
rect 149914 547574 150534 583018
rect 149914 547338 149946 547574
rect 150182 547338 150266 547574
rect 150502 547338 150534 547574
rect 149914 547254 150534 547338
rect 149914 547018 149946 547254
rect 150182 547018 150266 547254
rect 150502 547018 150534 547254
rect 149914 511574 150534 547018
rect 149914 511338 149946 511574
rect 150182 511338 150266 511574
rect 150502 511338 150534 511574
rect 149914 511254 150534 511338
rect 149914 511018 149946 511254
rect 150182 511018 150266 511254
rect 150502 511018 150534 511254
rect 149914 475574 150534 511018
rect 149914 475338 149946 475574
rect 150182 475338 150266 475574
rect 150502 475338 150534 475574
rect 149914 475254 150534 475338
rect 149914 475018 149946 475254
rect 150182 475018 150266 475254
rect 150502 475018 150534 475254
rect 149914 439574 150534 475018
rect 149914 439338 149946 439574
rect 150182 439338 150266 439574
rect 150502 439338 150534 439574
rect 149914 439254 150534 439338
rect 149914 439018 149946 439254
rect 150182 439018 150266 439254
rect 150502 439018 150534 439254
rect 149914 403574 150534 439018
rect 149914 403338 149946 403574
rect 150182 403338 150266 403574
rect 150502 403338 150534 403574
rect 149914 403254 150534 403338
rect 149914 403018 149946 403254
rect 150182 403018 150266 403254
rect 150502 403018 150534 403254
rect 149914 367574 150534 403018
rect 149914 367338 149946 367574
rect 150182 367338 150266 367574
rect 150502 367338 150534 367574
rect 149914 367254 150534 367338
rect 149914 367018 149946 367254
rect 150182 367018 150266 367254
rect 150502 367018 150534 367254
rect 149914 331574 150534 367018
rect 149914 331338 149946 331574
rect 150182 331338 150266 331574
rect 150502 331338 150534 331574
rect 149914 331254 150534 331338
rect 149914 331018 149946 331254
rect 150182 331018 150266 331254
rect 150502 331018 150534 331254
rect 149914 295574 150534 331018
rect 149914 295338 149946 295574
rect 150182 295338 150266 295574
rect 150502 295338 150534 295574
rect 149914 295254 150534 295338
rect 149914 295018 149946 295254
rect 150182 295018 150266 295254
rect 150502 295018 150534 295254
rect 149914 259574 150534 295018
rect 149914 259338 149946 259574
rect 150182 259338 150266 259574
rect 150502 259338 150534 259574
rect 149914 259254 150534 259338
rect 149914 259018 149946 259254
rect 150182 259018 150266 259254
rect 150502 259018 150534 259254
rect 149914 223574 150534 259018
rect 149914 223338 149946 223574
rect 150182 223338 150266 223574
rect 150502 223338 150534 223574
rect 149914 223254 150534 223338
rect 149914 223018 149946 223254
rect 150182 223018 150266 223254
rect 150502 223018 150534 223254
rect 149914 188457 150534 223018
rect 153634 706758 154254 711590
rect 153634 706522 153666 706758
rect 153902 706522 153986 706758
rect 154222 706522 154254 706758
rect 153634 706438 154254 706522
rect 153634 706202 153666 706438
rect 153902 706202 153986 706438
rect 154222 706202 154254 706438
rect 153634 695294 154254 706202
rect 153634 695058 153666 695294
rect 153902 695058 153986 695294
rect 154222 695058 154254 695294
rect 153634 694974 154254 695058
rect 153634 694738 153666 694974
rect 153902 694738 153986 694974
rect 154222 694738 154254 694974
rect 153634 659294 154254 694738
rect 153634 659058 153666 659294
rect 153902 659058 153986 659294
rect 154222 659058 154254 659294
rect 153634 658974 154254 659058
rect 153634 658738 153666 658974
rect 153902 658738 153986 658974
rect 154222 658738 154254 658974
rect 153634 623294 154254 658738
rect 153634 623058 153666 623294
rect 153902 623058 153986 623294
rect 154222 623058 154254 623294
rect 153634 622974 154254 623058
rect 153634 622738 153666 622974
rect 153902 622738 153986 622974
rect 154222 622738 154254 622974
rect 153634 587294 154254 622738
rect 153634 587058 153666 587294
rect 153902 587058 153986 587294
rect 154222 587058 154254 587294
rect 153634 586974 154254 587058
rect 153634 586738 153666 586974
rect 153902 586738 153986 586974
rect 154222 586738 154254 586974
rect 153634 551294 154254 586738
rect 153634 551058 153666 551294
rect 153902 551058 153986 551294
rect 154222 551058 154254 551294
rect 153634 550974 154254 551058
rect 153634 550738 153666 550974
rect 153902 550738 153986 550974
rect 154222 550738 154254 550974
rect 153634 515294 154254 550738
rect 153634 515058 153666 515294
rect 153902 515058 153986 515294
rect 154222 515058 154254 515294
rect 153634 514974 154254 515058
rect 153634 514738 153666 514974
rect 153902 514738 153986 514974
rect 154222 514738 154254 514974
rect 153634 479294 154254 514738
rect 153634 479058 153666 479294
rect 153902 479058 153986 479294
rect 154222 479058 154254 479294
rect 153634 478974 154254 479058
rect 153634 478738 153666 478974
rect 153902 478738 153986 478974
rect 154222 478738 154254 478974
rect 153634 443294 154254 478738
rect 153634 443058 153666 443294
rect 153902 443058 153986 443294
rect 154222 443058 154254 443294
rect 153634 442974 154254 443058
rect 153634 442738 153666 442974
rect 153902 442738 153986 442974
rect 154222 442738 154254 442974
rect 153634 407294 154254 442738
rect 153634 407058 153666 407294
rect 153902 407058 153986 407294
rect 154222 407058 154254 407294
rect 153634 406974 154254 407058
rect 153634 406738 153666 406974
rect 153902 406738 153986 406974
rect 154222 406738 154254 406974
rect 153634 371294 154254 406738
rect 153634 371058 153666 371294
rect 153902 371058 153986 371294
rect 154222 371058 154254 371294
rect 153634 370974 154254 371058
rect 153634 370738 153666 370974
rect 153902 370738 153986 370974
rect 154222 370738 154254 370974
rect 153634 335294 154254 370738
rect 153634 335058 153666 335294
rect 153902 335058 153986 335294
rect 154222 335058 154254 335294
rect 153634 334974 154254 335058
rect 153634 334738 153666 334974
rect 153902 334738 153986 334974
rect 154222 334738 154254 334974
rect 153634 299294 154254 334738
rect 153634 299058 153666 299294
rect 153902 299058 153986 299294
rect 154222 299058 154254 299294
rect 153634 298974 154254 299058
rect 153634 298738 153666 298974
rect 153902 298738 153986 298974
rect 154222 298738 154254 298974
rect 153634 263294 154254 298738
rect 153634 263058 153666 263294
rect 153902 263058 153986 263294
rect 154222 263058 154254 263294
rect 153634 262974 154254 263058
rect 153634 262738 153666 262974
rect 153902 262738 153986 262974
rect 154222 262738 154254 262974
rect 153634 227294 154254 262738
rect 153634 227058 153666 227294
rect 153902 227058 153986 227294
rect 154222 227058 154254 227294
rect 153634 226974 154254 227058
rect 153634 226738 153666 226974
rect 153902 226738 153986 226974
rect 154222 226738 154254 226974
rect 153634 191294 154254 226738
rect 153634 191058 153666 191294
rect 153902 191058 153986 191294
rect 154222 191058 154254 191294
rect 153634 190974 154254 191058
rect 153634 190738 153666 190974
rect 153902 190738 153986 190974
rect 154222 190738 154254 190974
rect 153634 188457 154254 190738
rect 157354 707718 157974 711590
rect 157354 707482 157386 707718
rect 157622 707482 157706 707718
rect 157942 707482 157974 707718
rect 157354 707398 157974 707482
rect 157354 707162 157386 707398
rect 157622 707162 157706 707398
rect 157942 707162 157974 707398
rect 157354 699014 157974 707162
rect 157354 698778 157386 699014
rect 157622 698778 157706 699014
rect 157942 698778 157974 699014
rect 157354 698694 157974 698778
rect 157354 698458 157386 698694
rect 157622 698458 157706 698694
rect 157942 698458 157974 698694
rect 157354 663014 157974 698458
rect 157354 662778 157386 663014
rect 157622 662778 157706 663014
rect 157942 662778 157974 663014
rect 157354 662694 157974 662778
rect 157354 662458 157386 662694
rect 157622 662458 157706 662694
rect 157942 662458 157974 662694
rect 157354 627014 157974 662458
rect 157354 626778 157386 627014
rect 157622 626778 157706 627014
rect 157942 626778 157974 627014
rect 157354 626694 157974 626778
rect 157354 626458 157386 626694
rect 157622 626458 157706 626694
rect 157942 626458 157974 626694
rect 157354 591014 157974 626458
rect 157354 590778 157386 591014
rect 157622 590778 157706 591014
rect 157942 590778 157974 591014
rect 157354 590694 157974 590778
rect 157354 590458 157386 590694
rect 157622 590458 157706 590694
rect 157942 590458 157974 590694
rect 157354 555014 157974 590458
rect 157354 554778 157386 555014
rect 157622 554778 157706 555014
rect 157942 554778 157974 555014
rect 157354 554694 157974 554778
rect 157354 554458 157386 554694
rect 157622 554458 157706 554694
rect 157942 554458 157974 554694
rect 157354 519014 157974 554458
rect 157354 518778 157386 519014
rect 157622 518778 157706 519014
rect 157942 518778 157974 519014
rect 157354 518694 157974 518778
rect 157354 518458 157386 518694
rect 157622 518458 157706 518694
rect 157942 518458 157974 518694
rect 157354 483014 157974 518458
rect 157354 482778 157386 483014
rect 157622 482778 157706 483014
rect 157942 482778 157974 483014
rect 157354 482694 157974 482778
rect 157354 482458 157386 482694
rect 157622 482458 157706 482694
rect 157942 482458 157974 482694
rect 157354 447014 157974 482458
rect 157354 446778 157386 447014
rect 157622 446778 157706 447014
rect 157942 446778 157974 447014
rect 157354 446694 157974 446778
rect 157354 446458 157386 446694
rect 157622 446458 157706 446694
rect 157942 446458 157974 446694
rect 157354 411014 157974 446458
rect 157354 410778 157386 411014
rect 157622 410778 157706 411014
rect 157942 410778 157974 411014
rect 157354 410694 157974 410778
rect 157354 410458 157386 410694
rect 157622 410458 157706 410694
rect 157942 410458 157974 410694
rect 157354 375014 157974 410458
rect 157354 374778 157386 375014
rect 157622 374778 157706 375014
rect 157942 374778 157974 375014
rect 157354 374694 157974 374778
rect 157354 374458 157386 374694
rect 157622 374458 157706 374694
rect 157942 374458 157974 374694
rect 157354 339014 157974 374458
rect 157354 338778 157386 339014
rect 157622 338778 157706 339014
rect 157942 338778 157974 339014
rect 157354 338694 157974 338778
rect 157354 338458 157386 338694
rect 157622 338458 157706 338694
rect 157942 338458 157974 338694
rect 157354 303014 157974 338458
rect 157354 302778 157386 303014
rect 157622 302778 157706 303014
rect 157942 302778 157974 303014
rect 157354 302694 157974 302778
rect 157354 302458 157386 302694
rect 157622 302458 157706 302694
rect 157942 302458 157974 302694
rect 157354 267014 157974 302458
rect 157354 266778 157386 267014
rect 157622 266778 157706 267014
rect 157942 266778 157974 267014
rect 157354 266694 157974 266778
rect 157354 266458 157386 266694
rect 157622 266458 157706 266694
rect 157942 266458 157974 266694
rect 157354 231014 157974 266458
rect 157354 230778 157386 231014
rect 157622 230778 157706 231014
rect 157942 230778 157974 231014
rect 157354 230694 157974 230778
rect 157354 230458 157386 230694
rect 157622 230458 157706 230694
rect 157942 230458 157974 230694
rect 157354 195014 157974 230458
rect 157354 194778 157386 195014
rect 157622 194778 157706 195014
rect 157942 194778 157974 195014
rect 157354 194694 157974 194778
rect 157354 194458 157386 194694
rect 157622 194458 157706 194694
rect 157942 194458 157974 194694
rect 157354 188457 157974 194458
rect 161074 708678 161694 711590
rect 161074 708442 161106 708678
rect 161342 708442 161426 708678
rect 161662 708442 161694 708678
rect 161074 708358 161694 708442
rect 161074 708122 161106 708358
rect 161342 708122 161426 708358
rect 161662 708122 161694 708358
rect 161074 666734 161694 708122
rect 161074 666498 161106 666734
rect 161342 666498 161426 666734
rect 161662 666498 161694 666734
rect 161074 666414 161694 666498
rect 161074 666178 161106 666414
rect 161342 666178 161426 666414
rect 161662 666178 161694 666414
rect 161074 630734 161694 666178
rect 161074 630498 161106 630734
rect 161342 630498 161426 630734
rect 161662 630498 161694 630734
rect 161074 630414 161694 630498
rect 161074 630178 161106 630414
rect 161342 630178 161426 630414
rect 161662 630178 161694 630414
rect 161074 594734 161694 630178
rect 161074 594498 161106 594734
rect 161342 594498 161426 594734
rect 161662 594498 161694 594734
rect 161074 594414 161694 594498
rect 161074 594178 161106 594414
rect 161342 594178 161426 594414
rect 161662 594178 161694 594414
rect 161074 558734 161694 594178
rect 161074 558498 161106 558734
rect 161342 558498 161426 558734
rect 161662 558498 161694 558734
rect 161074 558414 161694 558498
rect 161074 558178 161106 558414
rect 161342 558178 161426 558414
rect 161662 558178 161694 558414
rect 161074 522734 161694 558178
rect 161074 522498 161106 522734
rect 161342 522498 161426 522734
rect 161662 522498 161694 522734
rect 161074 522414 161694 522498
rect 161074 522178 161106 522414
rect 161342 522178 161426 522414
rect 161662 522178 161694 522414
rect 161074 486734 161694 522178
rect 161074 486498 161106 486734
rect 161342 486498 161426 486734
rect 161662 486498 161694 486734
rect 161074 486414 161694 486498
rect 161074 486178 161106 486414
rect 161342 486178 161426 486414
rect 161662 486178 161694 486414
rect 161074 450734 161694 486178
rect 161074 450498 161106 450734
rect 161342 450498 161426 450734
rect 161662 450498 161694 450734
rect 161074 450414 161694 450498
rect 161074 450178 161106 450414
rect 161342 450178 161426 450414
rect 161662 450178 161694 450414
rect 161074 414734 161694 450178
rect 161074 414498 161106 414734
rect 161342 414498 161426 414734
rect 161662 414498 161694 414734
rect 161074 414414 161694 414498
rect 161074 414178 161106 414414
rect 161342 414178 161426 414414
rect 161662 414178 161694 414414
rect 161074 378734 161694 414178
rect 161074 378498 161106 378734
rect 161342 378498 161426 378734
rect 161662 378498 161694 378734
rect 161074 378414 161694 378498
rect 161074 378178 161106 378414
rect 161342 378178 161426 378414
rect 161662 378178 161694 378414
rect 161074 342734 161694 378178
rect 161074 342498 161106 342734
rect 161342 342498 161426 342734
rect 161662 342498 161694 342734
rect 161074 342414 161694 342498
rect 161074 342178 161106 342414
rect 161342 342178 161426 342414
rect 161662 342178 161694 342414
rect 161074 306734 161694 342178
rect 161074 306498 161106 306734
rect 161342 306498 161426 306734
rect 161662 306498 161694 306734
rect 161074 306414 161694 306498
rect 161074 306178 161106 306414
rect 161342 306178 161426 306414
rect 161662 306178 161694 306414
rect 161074 270734 161694 306178
rect 161074 270498 161106 270734
rect 161342 270498 161426 270734
rect 161662 270498 161694 270734
rect 161074 270414 161694 270498
rect 161074 270178 161106 270414
rect 161342 270178 161426 270414
rect 161662 270178 161694 270414
rect 161074 234734 161694 270178
rect 161074 234498 161106 234734
rect 161342 234498 161426 234734
rect 161662 234498 161694 234734
rect 161074 234414 161694 234498
rect 161074 234178 161106 234414
rect 161342 234178 161426 234414
rect 161662 234178 161694 234414
rect 161074 198734 161694 234178
rect 161074 198498 161106 198734
rect 161342 198498 161426 198734
rect 161662 198498 161694 198734
rect 161074 198414 161694 198498
rect 161074 198178 161106 198414
rect 161342 198178 161426 198414
rect 161662 198178 161694 198414
rect 161074 189900 161694 198178
rect 164794 709638 165414 711590
rect 164794 709402 164826 709638
rect 165062 709402 165146 709638
rect 165382 709402 165414 709638
rect 164794 709318 165414 709402
rect 164794 709082 164826 709318
rect 165062 709082 165146 709318
rect 165382 709082 165414 709318
rect 164794 670454 165414 709082
rect 164794 670218 164826 670454
rect 165062 670218 165146 670454
rect 165382 670218 165414 670454
rect 164794 670134 165414 670218
rect 164794 669898 164826 670134
rect 165062 669898 165146 670134
rect 165382 669898 165414 670134
rect 164794 634454 165414 669898
rect 164794 634218 164826 634454
rect 165062 634218 165146 634454
rect 165382 634218 165414 634454
rect 164794 634134 165414 634218
rect 164794 633898 164826 634134
rect 165062 633898 165146 634134
rect 165382 633898 165414 634134
rect 164794 598454 165414 633898
rect 164794 598218 164826 598454
rect 165062 598218 165146 598454
rect 165382 598218 165414 598454
rect 164794 598134 165414 598218
rect 164794 597898 164826 598134
rect 165062 597898 165146 598134
rect 165382 597898 165414 598134
rect 164794 562454 165414 597898
rect 164794 562218 164826 562454
rect 165062 562218 165146 562454
rect 165382 562218 165414 562454
rect 164794 562134 165414 562218
rect 164794 561898 164826 562134
rect 165062 561898 165146 562134
rect 165382 561898 165414 562134
rect 164794 526454 165414 561898
rect 164794 526218 164826 526454
rect 165062 526218 165146 526454
rect 165382 526218 165414 526454
rect 164794 526134 165414 526218
rect 164794 525898 164826 526134
rect 165062 525898 165146 526134
rect 165382 525898 165414 526134
rect 164794 490454 165414 525898
rect 164794 490218 164826 490454
rect 165062 490218 165146 490454
rect 165382 490218 165414 490454
rect 164794 490134 165414 490218
rect 164794 489898 164826 490134
rect 165062 489898 165146 490134
rect 165382 489898 165414 490134
rect 164794 454454 165414 489898
rect 164794 454218 164826 454454
rect 165062 454218 165146 454454
rect 165382 454218 165414 454454
rect 164794 454134 165414 454218
rect 164794 453898 164826 454134
rect 165062 453898 165146 454134
rect 165382 453898 165414 454134
rect 164794 418454 165414 453898
rect 164794 418218 164826 418454
rect 165062 418218 165146 418454
rect 165382 418218 165414 418454
rect 164794 418134 165414 418218
rect 164794 417898 164826 418134
rect 165062 417898 165146 418134
rect 165382 417898 165414 418134
rect 164794 382454 165414 417898
rect 164794 382218 164826 382454
rect 165062 382218 165146 382454
rect 165382 382218 165414 382454
rect 164794 382134 165414 382218
rect 164794 381898 164826 382134
rect 165062 381898 165146 382134
rect 165382 381898 165414 382134
rect 164794 346454 165414 381898
rect 164794 346218 164826 346454
rect 165062 346218 165146 346454
rect 165382 346218 165414 346454
rect 164794 346134 165414 346218
rect 164794 345898 164826 346134
rect 165062 345898 165146 346134
rect 165382 345898 165414 346134
rect 164794 310454 165414 345898
rect 164794 310218 164826 310454
rect 165062 310218 165146 310454
rect 165382 310218 165414 310454
rect 164794 310134 165414 310218
rect 164794 309898 164826 310134
rect 165062 309898 165146 310134
rect 165382 309898 165414 310134
rect 164794 274454 165414 309898
rect 164794 274218 164826 274454
rect 165062 274218 165146 274454
rect 165382 274218 165414 274454
rect 164794 274134 165414 274218
rect 164794 273898 164826 274134
rect 165062 273898 165146 274134
rect 165382 273898 165414 274134
rect 164794 238454 165414 273898
rect 164794 238218 164826 238454
rect 165062 238218 165146 238454
rect 165382 238218 165414 238454
rect 164794 238134 165414 238218
rect 164794 237898 164826 238134
rect 165062 237898 165146 238134
rect 165382 237898 165414 238134
rect 164794 202454 165414 237898
rect 164794 202218 164826 202454
rect 165062 202218 165146 202454
rect 165382 202218 165414 202454
rect 164794 202134 165414 202218
rect 164794 201898 164826 202134
rect 165062 201898 165146 202134
rect 165382 201898 165414 202134
rect 164794 188457 165414 201898
rect 168514 710598 169134 711590
rect 168514 710362 168546 710598
rect 168782 710362 168866 710598
rect 169102 710362 169134 710598
rect 168514 710278 169134 710362
rect 168514 710042 168546 710278
rect 168782 710042 168866 710278
rect 169102 710042 169134 710278
rect 168514 674174 169134 710042
rect 168514 673938 168546 674174
rect 168782 673938 168866 674174
rect 169102 673938 169134 674174
rect 168514 673854 169134 673938
rect 168514 673618 168546 673854
rect 168782 673618 168866 673854
rect 169102 673618 169134 673854
rect 168514 638174 169134 673618
rect 168514 637938 168546 638174
rect 168782 637938 168866 638174
rect 169102 637938 169134 638174
rect 168514 637854 169134 637938
rect 168514 637618 168546 637854
rect 168782 637618 168866 637854
rect 169102 637618 169134 637854
rect 168514 602174 169134 637618
rect 168514 601938 168546 602174
rect 168782 601938 168866 602174
rect 169102 601938 169134 602174
rect 168514 601854 169134 601938
rect 168514 601618 168546 601854
rect 168782 601618 168866 601854
rect 169102 601618 169134 601854
rect 168514 566174 169134 601618
rect 168514 565938 168546 566174
rect 168782 565938 168866 566174
rect 169102 565938 169134 566174
rect 168514 565854 169134 565938
rect 168514 565618 168546 565854
rect 168782 565618 168866 565854
rect 169102 565618 169134 565854
rect 168514 530174 169134 565618
rect 168514 529938 168546 530174
rect 168782 529938 168866 530174
rect 169102 529938 169134 530174
rect 168514 529854 169134 529938
rect 168514 529618 168546 529854
rect 168782 529618 168866 529854
rect 169102 529618 169134 529854
rect 168514 494174 169134 529618
rect 168514 493938 168546 494174
rect 168782 493938 168866 494174
rect 169102 493938 169134 494174
rect 168514 493854 169134 493938
rect 168514 493618 168546 493854
rect 168782 493618 168866 493854
rect 169102 493618 169134 493854
rect 168514 458174 169134 493618
rect 168514 457938 168546 458174
rect 168782 457938 168866 458174
rect 169102 457938 169134 458174
rect 168514 457854 169134 457938
rect 168514 457618 168546 457854
rect 168782 457618 168866 457854
rect 169102 457618 169134 457854
rect 168514 422174 169134 457618
rect 168514 421938 168546 422174
rect 168782 421938 168866 422174
rect 169102 421938 169134 422174
rect 168514 421854 169134 421938
rect 168514 421618 168546 421854
rect 168782 421618 168866 421854
rect 169102 421618 169134 421854
rect 168514 386174 169134 421618
rect 168514 385938 168546 386174
rect 168782 385938 168866 386174
rect 169102 385938 169134 386174
rect 168514 385854 169134 385938
rect 168514 385618 168546 385854
rect 168782 385618 168866 385854
rect 169102 385618 169134 385854
rect 168514 350174 169134 385618
rect 168514 349938 168546 350174
rect 168782 349938 168866 350174
rect 169102 349938 169134 350174
rect 168514 349854 169134 349938
rect 168514 349618 168546 349854
rect 168782 349618 168866 349854
rect 169102 349618 169134 349854
rect 168514 314174 169134 349618
rect 168514 313938 168546 314174
rect 168782 313938 168866 314174
rect 169102 313938 169134 314174
rect 168514 313854 169134 313938
rect 168514 313618 168546 313854
rect 168782 313618 168866 313854
rect 169102 313618 169134 313854
rect 168514 278174 169134 313618
rect 168514 277938 168546 278174
rect 168782 277938 168866 278174
rect 169102 277938 169134 278174
rect 168514 277854 169134 277938
rect 168514 277618 168546 277854
rect 168782 277618 168866 277854
rect 169102 277618 169134 277854
rect 168514 242174 169134 277618
rect 168514 241938 168546 242174
rect 168782 241938 168866 242174
rect 169102 241938 169134 242174
rect 168514 241854 169134 241938
rect 168514 241618 168546 241854
rect 168782 241618 168866 241854
rect 169102 241618 169134 241854
rect 168514 206174 169134 241618
rect 168514 205938 168546 206174
rect 168782 205938 168866 206174
rect 169102 205938 169134 206174
rect 168514 205854 169134 205938
rect 168514 205618 168546 205854
rect 168782 205618 168866 205854
rect 169102 205618 169134 205854
rect 168514 188457 169134 205618
rect 172234 711558 172854 711590
rect 172234 711322 172266 711558
rect 172502 711322 172586 711558
rect 172822 711322 172854 711558
rect 172234 711238 172854 711322
rect 172234 711002 172266 711238
rect 172502 711002 172586 711238
rect 172822 711002 172854 711238
rect 172234 677894 172854 711002
rect 172234 677658 172266 677894
rect 172502 677658 172586 677894
rect 172822 677658 172854 677894
rect 172234 677574 172854 677658
rect 172234 677338 172266 677574
rect 172502 677338 172586 677574
rect 172822 677338 172854 677574
rect 172234 641894 172854 677338
rect 172234 641658 172266 641894
rect 172502 641658 172586 641894
rect 172822 641658 172854 641894
rect 172234 641574 172854 641658
rect 172234 641338 172266 641574
rect 172502 641338 172586 641574
rect 172822 641338 172854 641574
rect 172234 605894 172854 641338
rect 172234 605658 172266 605894
rect 172502 605658 172586 605894
rect 172822 605658 172854 605894
rect 172234 605574 172854 605658
rect 172234 605338 172266 605574
rect 172502 605338 172586 605574
rect 172822 605338 172854 605574
rect 172234 569894 172854 605338
rect 172234 569658 172266 569894
rect 172502 569658 172586 569894
rect 172822 569658 172854 569894
rect 172234 569574 172854 569658
rect 172234 569338 172266 569574
rect 172502 569338 172586 569574
rect 172822 569338 172854 569574
rect 172234 533894 172854 569338
rect 172234 533658 172266 533894
rect 172502 533658 172586 533894
rect 172822 533658 172854 533894
rect 172234 533574 172854 533658
rect 172234 533338 172266 533574
rect 172502 533338 172586 533574
rect 172822 533338 172854 533574
rect 172234 497894 172854 533338
rect 172234 497658 172266 497894
rect 172502 497658 172586 497894
rect 172822 497658 172854 497894
rect 172234 497574 172854 497658
rect 172234 497338 172266 497574
rect 172502 497338 172586 497574
rect 172822 497338 172854 497574
rect 172234 461894 172854 497338
rect 172234 461658 172266 461894
rect 172502 461658 172586 461894
rect 172822 461658 172854 461894
rect 172234 461574 172854 461658
rect 172234 461338 172266 461574
rect 172502 461338 172586 461574
rect 172822 461338 172854 461574
rect 172234 425894 172854 461338
rect 172234 425658 172266 425894
rect 172502 425658 172586 425894
rect 172822 425658 172854 425894
rect 172234 425574 172854 425658
rect 172234 425338 172266 425574
rect 172502 425338 172586 425574
rect 172822 425338 172854 425574
rect 172234 389894 172854 425338
rect 172234 389658 172266 389894
rect 172502 389658 172586 389894
rect 172822 389658 172854 389894
rect 172234 389574 172854 389658
rect 172234 389338 172266 389574
rect 172502 389338 172586 389574
rect 172822 389338 172854 389574
rect 172234 353894 172854 389338
rect 172234 353658 172266 353894
rect 172502 353658 172586 353894
rect 172822 353658 172854 353894
rect 172234 353574 172854 353658
rect 172234 353338 172266 353574
rect 172502 353338 172586 353574
rect 172822 353338 172854 353574
rect 172234 317894 172854 353338
rect 172234 317658 172266 317894
rect 172502 317658 172586 317894
rect 172822 317658 172854 317894
rect 172234 317574 172854 317658
rect 172234 317338 172266 317574
rect 172502 317338 172586 317574
rect 172822 317338 172854 317574
rect 172234 281894 172854 317338
rect 172234 281658 172266 281894
rect 172502 281658 172586 281894
rect 172822 281658 172854 281894
rect 172234 281574 172854 281658
rect 172234 281338 172266 281574
rect 172502 281338 172586 281574
rect 172822 281338 172854 281574
rect 172234 245894 172854 281338
rect 172234 245658 172266 245894
rect 172502 245658 172586 245894
rect 172822 245658 172854 245894
rect 172234 245574 172854 245658
rect 172234 245338 172266 245574
rect 172502 245338 172586 245574
rect 172822 245338 172854 245574
rect 172234 209894 172854 245338
rect 172234 209658 172266 209894
rect 172502 209658 172586 209894
rect 172822 209658 172854 209894
rect 172234 209574 172854 209658
rect 172234 209338 172266 209574
rect 172502 209338 172586 209574
rect 172822 209338 172854 209574
rect 172234 188457 172854 209338
rect 182194 704838 182814 711590
rect 182194 704602 182226 704838
rect 182462 704602 182546 704838
rect 182782 704602 182814 704838
rect 182194 704518 182814 704602
rect 182194 704282 182226 704518
rect 182462 704282 182546 704518
rect 182782 704282 182814 704518
rect 182194 687854 182814 704282
rect 182194 687618 182226 687854
rect 182462 687618 182546 687854
rect 182782 687618 182814 687854
rect 182194 687534 182814 687618
rect 182194 687298 182226 687534
rect 182462 687298 182546 687534
rect 182782 687298 182814 687534
rect 182194 651854 182814 687298
rect 182194 651618 182226 651854
rect 182462 651618 182546 651854
rect 182782 651618 182814 651854
rect 182194 651534 182814 651618
rect 182194 651298 182226 651534
rect 182462 651298 182546 651534
rect 182782 651298 182814 651534
rect 182194 615854 182814 651298
rect 182194 615618 182226 615854
rect 182462 615618 182546 615854
rect 182782 615618 182814 615854
rect 182194 615534 182814 615618
rect 182194 615298 182226 615534
rect 182462 615298 182546 615534
rect 182782 615298 182814 615534
rect 182194 579854 182814 615298
rect 182194 579618 182226 579854
rect 182462 579618 182546 579854
rect 182782 579618 182814 579854
rect 182194 579534 182814 579618
rect 182194 579298 182226 579534
rect 182462 579298 182546 579534
rect 182782 579298 182814 579534
rect 182194 543854 182814 579298
rect 182194 543618 182226 543854
rect 182462 543618 182546 543854
rect 182782 543618 182814 543854
rect 182194 543534 182814 543618
rect 182194 543298 182226 543534
rect 182462 543298 182546 543534
rect 182782 543298 182814 543534
rect 182194 507854 182814 543298
rect 182194 507618 182226 507854
rect 182462 507618 182546 507854
rect 182782 507618 182814 507854
rect 182194 507534 182814 507618
rect 182194 507298 182226 507534
rect 182462 507298 182546 507534
rect 182782 507298 182814 507534
rect 182194 471854 182814 507298
rect 182194 471618 182226 471854
rect 182462 471618 182546 471854
rect 182782 471618 182814 471854
rect 182194 471534 182814 471618
rect 182194 471298 182226 471534
rect 182462 471298 182546 471534
rect 182782 471298 182814 471534
rect 182194 435854 182814 471298
rect 182194 435618 182226 435854
rect 182462 435618 182546 435854
rect 182782 435618 182814 435854
rect 182194 435534 182814 435618
rect 182194 435298 182226 435534
rect 182462 435298 182546 435534
rect 182782 435298 182814 435534
rect 182194 399854 182814 435298
rect 182194 399618 182226 399854
rect 182462 399618 182546 399854
rect 182782 399618 182814 399854
rect 182194 399534 182814 399618
rect 182194 399298 182226 399534
rect 182462 399298 182546 399534
rect 182782 399298 182814 399534
rect 182194 363854 182814 399298
rect 182194 363618 182226 363854
rect 182462 363618 182546 363854
rect 182782 363618 182814 363854
rect 182194 363534 182814 363618
rect 182194 363298 182226 363534
rect 182462 363298 182546 363534
rect 182782 363298 182814 363534
rect 182194 327854 182814 363298
rect 182194 327618 182226 327854
rect 182462 327618 182546 327854
rect 182782 327618 182814 327854
rect 182194 327534 182814 327618
rect 182194 327298 182226 327534
rect 182462 327298 182546 327534
rect 182782 327298 182814 327534
rect 182194 291854 182814 327298
rect 182194 291618 182226 291854
rect 182462 291618 182546 291854
rect 182782 291618 182814 291854
rect 182194 291534 182814 291618
rect 182194 291298 182226 291534
rect 182462 291298 182546 291534
rect 182782 291298 182814 291534
rect 182194 255854 182814 291298
rect 182194 255618 182226 255854
rect 182462 255618 182546 255854
rect 182782 255618 182814 255854
rect 182194 255534 182814 255618
rect 182194 255298 182226 255534
rect 182462 255298 182546 255534
rect 182782 255298 182814 255534
rect 182194 219854 182814 255298
rect 182194 219618 182226 219854
rect 182462 219618 182546 219854
rect 182782 219618 182814 219854
rect 182194 219534 182814 219618
rect 182194 219298 182226 219534
rect 182462 219298 182546 219534
rect 182782 219298 182814 219534
rect 182194 188457 182814 219298
rect 185914 705798 186534 711590
rect 185914 705562 185946 705798
rect 186182 705562 186266 705798
rect 186502 705562 186534 705798
rect 185914 705478 186534 705562
rect 185914 705242 185946 705478
rect 186182 705242 186266 705478
rect 186502 705242 186534 705478
rect 185914 691574 186534 705242
rect 185914 691338 185946 691574
rect 186182 691338 186266 691574
rect 186502 691338 186534 691574
rect 185914 691254 186534 691338
rect 185914 691018 185946 691254
rect 186182 691018 186266 691254
rect 186502 691018 186534 691254
rect 185914 655574 186534 691018
rect 185914 655338 185946 655574
rect 186182 655338 186266 655574
rect 186502 655338 186534 655574
rect 185914 655254 186534 655338
rect 185914 655018 185946 655254
rect 186182 655018 186266 655254
rect 186502 655018 186534 655254
rect 185914 619574 186534 655018
rect 185914 619338 185946 619574
rect 186182 619338 186266 619574
rect 186502 619338 186534 619574
rect 185914 619254 186534 619338
rect 185914 619018 185946 619254
rect 186182 619018 186266 619254
rect 186502 619018 186534 619254
rect 185914 583574 186534 619018
rect 185914 583338 185946 583574
rect 186182 583338 186266 583574
rect 186502 583338 186534 583574
rect 185914 583254 186534 583338
rect 185914 583018 185946 583254
rect 186182 583018 186266 583254
rect 186502 583018 186534 583254
rect 185914 547574 186534 583018
rect 185914 547338 185946 547574
rect 186182 547338 186266 547574
rect 186502 547338 186534 547574
rect 185914 547254 186534 547338
rect 185914 547018 185946 547254
rect 186182 547018 186266 547254
rect 186502 547018 186534 547254
rect 185914 511574 186534 547018
rect 185914 511338 185946 511574
rect 186182 511338 186266 511574
rect 186502 511338 186534 511574
rect 185914 511254 186534 511338
rect 185914 511018 185946 511254
rect 186182 511018 186266 511254
rect 186502 511018 186534 511254
rect 185914 475574 186534 511018
rect 185914 475338 185946 475574
rect 186182 475338 186266 475574
rect 186502 475338 186534 475574
rect 185914 475254 186534 475338
rect 185914 475018 185946 475254
rect 186182 475018 186266 475254
rect 186502 475018 186534 475254
rect 185914 439574 186534 475018
rect 185914 439338 185946 439574
rect 186182 439338 186266 439574
rect 186502 439338 186534 439574
rect 185914 439254 186534 439338
rect 185914 439018 185946 439254
rect 186182 439018 186266 439254
rect 186502 439018 186534 439254
rect 185914 403574 186534 439018
rect 185914 403338 185946 403574
rect 186182 403338 186266 403574
rect 186502 403338 186534 403574
rect 185914 403254 186534 403338
rect 185914 403018 185946 403254
rect 186182 403018 186266 403254
rect 186502 403018 186534 403254
rect 185914 367574 186534 403018
rect 185914 367338 185946 367574
rect 186182 367338 186266 367574
rect 186502 367338 186534 367574
rect 185914 367254 186534 367338
rect 185914 367018 185946 367254
rect 186182 367018 186266 367254
rect 186502 367018 186534 367254
rect 185914 331574 186534 367018
rect 185914 331338 185946 331574
rect 186182 331338 186266 331574
rect 186502 331338 186534 331574
rect 185914 331254 186534 331338
rect 185914 331018 185946 331254
rect 186182 331018 186266 331254
rect 186502 331018 186534 331254
rect 185914 295574 186534 331018
rect 185914 295338 185946 295574
rect 186182 295338 186266 295574
rect 186502 295338 186534 295574
rect 185914 295254 186534 295338
rect 185914 295018 185946 295254
rect 186182 295018 186266 295254
rect 186502 295018 186534 295254
rect 185914 259574 186534 295018
rect 185914 259338 185946 259574
rect 186182 259338 186266 259574
rect 186502 259338 186534 259574
rect 185914 259254 186534 259338
rect 185914 259018 185946 259254
rect 186182 259018 186266 259254
rect 186502 259018 186534 259254
rect 185914 223574 186534 259018
rect 185914 223338 185946 223574
rect 186182 223338 186266 223574
rect 186502 223338 186534 223574
rect 185914 223254 186534 223338
rect 185914 223018 185946 223254
rect 186182 223018 186266 223254
rect 186502 223018 186534 223254
rect 185914 188457 186534 223018
rect 189634 706758 190254 711590
rect 189634 706522 189666 706758
rect 189902 706522 189986 706758
rect 190222 706522 190254 706758
rect 189634 706438 190254 706522
rect 189634 706202 189666 706438
rect 189902 706202 189986 706438
rect 190222 706202 190254 706438
rect 189634 695294 190254 706202
rect 193354 707718 193974 711590
rect 193354 707482 193386 707718
rect 193622 707482 193706 707718
rect 193942 707482 193974 707718
rect 193354 707398 193974 707482
rect 193354 707162 193386 707398
rect 193622 707162 193706 707398
rect 193942 707162 193974 707398
rect 192339 700500 192405 700501
rect 192339 700436 192340 700500
rect 192404 700436 192405 700500
rect 192339 700435 192405 700436
rect 189634 695058 189666 695294
rect 189902 695058 189986 695294
rect 190222 695058 190254 695294
rect 189634 694974 190254 695058
rect 189634 694738 189666 694974
rect 189902 694738 189986 694974
rect 190222 694738 190254 694974
rect 189634 659294 190254 694738
rect 189634 659058 189666 659294
rect 189902 659058 189986 659294
rect 190222 659058 190254 659294
rect 189634 658974 190254 659058
rect 189634 658738 189666 658974
rect 189902 658738 189986 658974
rect 190222 658738 190254 658974
rect 189634 623294 190254 658738
rect 189634 623058 189666 623294
rect 189902 623058 189986 623294
rect 190222 623058 190254 623294
rect 189634 622974 190254 623058
rect 189634 622738 189666 622974
rect 189902 622738 189986 622974
rect 190222 622738 190254 622974
rect 189634 587294 190254 622738
rect 189634 587058 189666 587294
rect 189902 587058 189986 587294
rect 190222 587058 190254 587294
rect 189634 586974 190254 587058
rect 189634 586738 189666 586974
rect 189902 586738 189986 586974
rect 190222 586738 190254 586974
rect 189634 551294 190254 586738
rect 189634 551058 189666 551294
rect 189902 551058 189986 551294
rect 190222 551058 190254 551294
rect 189634 550974 190254 551058
rect 189634 550738 189666 550974
rect 189902 550738 189986 550974
rect 190222 550738 190254 550974
rect 189634 515294 190254 550738
rect 189634 515058 189666 515294
rect 189902 515058 189986 515294
rect 190222 515058 190254 515294
rect 189634 514974 190254 515058
rect 189634 514738 189666 514974
rect 189902 514738 189986 514974
rect 190222 514738 190254 514974
rect 189634 479294 190254 514738
rect 189634 479058 189666 479294
rect 189902 479058 189986 479294
rect 190222 479058 190254 479294
rect 189634 478974 190254 479058
rect 189634 478738 189666 478974
rect 189902 478738 189986 478974
rect 190222 478738 190254 478974
rect 189634 443294 190254 478738
rect 189634 443058 189666 443294
rect 189902 443058 189986 443294
rect 190222 443058 190254 443294
rect 189634 442974 190254 443058
rect 189634 442738 189666 442974
rect 189902 442738 189986 442974
rect 190222 442738 190254 442974
rect 189634 407294 190254 442738
rect 189634 407058 189666 407294
rect 189902 407058 189986 407294
rect 190222 407058 190254 407294
rect 189634 406974 190254 407058
rect 189634 406738 189666 406974
rect 189902 406738 189986 406974
rect 190222 406738 190254 406974
rect 189634 371294 190254 406738
rect 189634 371058 189666 371294
rect 189902 371058 189986 371294
rect 190222 371058 190254 371294
rect 189634 370974 190254 371058
rect 189634 370738 189666 370974
rect 189902 370738 189986 370974
rect 190222 370738 190254 370974
rect 189634 335294 190254 370738
rect 189634 335058 189666 335294
rect 189902 335058 189986 335294
rect 190222 335058 190254 335294
rect 189634 334974 190254 335058
rect 189634 334738 189666 334974
rect 189902 334738 189986 334974
rect 190222 334738 190254 334974
rect 189634 299294 190254 334738
rect 189634 299058 189666 299294
rect 189902 299058 189986 299294
rect 190222 299058 190254 299294
rect 189634 298974 190254 299058
rect 189634 298738 189666 298974
rect 189902 298738 189986 298974
rect 190222 298738 190254 298974
rect 189634 263294 190254 298738
rect 189634 263058 189666 263294
rect 189902 263058 189986 263294
rect 190222 263058 190254 263294
rect 189634 262974 190254 263058
rect 189634 262738 189666 262974
rect 189902 262738 189986 262974
rect 190222 262738 190254 262974
rect 189634 227294 190254 262738
rect 189634 227058 189666 227294
rect 189902 227058 189986 227294
rect 190222 227058 190254 227294
rect 189634 226974 190254 227058
rect 189634 226738 189666 226974
rect 189902 226738 189986 226974
rect 190222 226738 190254 226974
rect 189634 191294 190254 226738
rect 189634 191058 189666 191294
rect 189902 191058 189986 191294
rect 190222 191058 190254 191294
rect 189634 190974 190254 191058
rect 189634 190738 189666 190974
rect 189902 190738 189986 190974
rect 190222 190738 190254 190974
rect 99568 187574 99888 187606
rect 99568 187338 99610 187574
rect 99846 187338 99888 187574
rect 99568 187254 99888 187338
rect 99568 187018 99610 187254
rect 99846 187018 99888 187254
rect 99568 186986 99888 187018
rect 130288 187574 130608 187606
rect 130288 187338 130330 187574
rect 130566 187338 130608 187574
rect 130288 187254 130608 187338
rect 130288 187018 130330 187254
rect 130566 187018 130608 187254
rect 130288 186986 130608 187018
rect 161008 187574 161328 187606
rect 161008 187338 161050 187574
rect 161286 187338 161328 187574
rect 161008 187254 161328 187338
rect 161008 187018 161050 187254
rect 161286 187018 161328 187254
rect 161008 186986 161328 187018
rect 114928 183854 115248 183886
rect 114928 183618 114970 183854
rect 115206 183618 115248 183854
rect 114928 183534 115248 183618
rect 114928 183298 114970 183534
rect 115206 183298 115248 183534
rect 114928 183266 115248 183298
rect 145648 183854 145968 183886
rect 145648 183618 145690 183854
rect 145926 183618 145968 183854
rect 145648 183534 145968 183618
rect 145648 183298 145690 183534
rect 145926 183298 145968 183534
rect 145648 183266 145968 183298
rect 176368 183854 176688 183886
rect 176368 183618 176410 183854
rect 176646 183618 176688 183854
rect 176368 183534 176688 183618
rect 176368 183298 176410 183534
rect 176646 183298 176688 183534
rect 176368 183266 176688 183298
rect 96514 169938 96546 170174
rect 96782 169938 96866 170174
rect 97102 169938 97134 170174
rect 96514 169854 97134 169938
rect 96514 169618 96546 169854
rect 96782 169618 96866 169854
rect 97102 169618 97134 169854
rect 96514 134174 97134 169618
rect 189634 155294 190254 190738
rect 191787 177172 191853 177173
rect 191787 177108 191788 177172
rect 191852 177108 191853 177172
rect 191787 177107 191853 177108
rect 189634 155058 189666 155294
rect 189902 155058 189986 155294
rect 190222 155058 190254 155294
rect 189634 154974 190254 155058
rect 189634 154738 189666 154974
rect 189902 154738 189986 154974
rect 190222 154738 190254 154974
rect 99568 151574 99888 151606
rect 99568 151338 99610 151574
rect 99846 151338 99888 151574
rect 99568 151254 99888 151338
rect 99568 151018 99610 151254
rect 99846 151018 99888 151254
rect 99568 150986 99888 151018
rect 130288 151574 130608 151606
rect 130288 151338 130330 151574
rect 130566 151338 130608 151574
rect 130288 151254 130608 151338
rect 130288 151018 130330 151254
rect 130566 151018 130608 151254
rect 130288 150986 130608 151018
rect 161008 151574 161328 151606
rect 161008 151338 161050 151574
rect 161286 151338 161328 151574
rect 161008 151254 161328 151338
rect 161008 151018 161050 151254
rect 161286 151018 161328 151254
rect 161008 150986 161328 151018
rect 114928 147854 115248 147886
rect 114928 147618 114970 147854
rect 115206 147618 115248 147854
rect 114928 147534 115248 147618
rect 114928 147298 114970 147534
rect 115206 147298 115248 147534
rect 114928 147266 115248 147298
rect 145648 147854 145968 147886
rect 145648 147618 145690 147854
rect 145926 147618 145968 147854
rect 145648 147534 145968 147618
rect 145648 147298 145690 147534
rect 145926 147298 145968 147534
rect 145648 147266 145968 147298
rect 176368 147854 176688 147886
rect 176368 147618 176410 147854
rect 176646 147618 176688 147854
rect 176368 147534 176688 147618
rect 176368 147298 176410 147534
rect 176646 147298 176688 147534
rect 176368 147266 176688 147298
rect 96514 133938 96546 134174
rect 96782 133938 96866 134174
rect 97102 133938 97134 134174
rect 96514 133854 97134 133938
rect 96514 133618 96546 133854
rect 96782 133618 96866 133854
rect 97102 133618 97134 133854
rect 96514 98174 97134 133618
rect 189634 119294 190254 154738
rect 191235 127124 191301 127125
rect 191235 127060 191236 127124
rect 191300 127060 191301 127124
rect 191235 127059 191301 127060
rect 189634 119058 189666 119294
rect 189902 119058 189986 119294
rect 190222 119058 190254 119294
rect 189634 118974 190254 119058
rect 189634 118738 189666 118974
rect 189902 118738 189986 118974
rect 190222 118738 190254 118974
rect 99568 115574 99888 115606
rect 99568 115338 99610 115574
rect 99846 115338 99888 115574
rect 99568 115254 99888 115338
rect 99568 115018 99610 115254
rect 99846 115018 99888 115254
rect 99568 114986 99888 115018
rect 130288 115574 130608 115606
rect 130288 115338 130330 115574
rect 130566 115338 130608 115574
rect 130288 115254 130608 115338
rect 130288 115018 130330 115254
rect 130566 115018 130608 115254
rect 130288 114986 130608 115018
rect 161008 115574 161328 115606
rect 161008 115338 161050 115574
rect 161286 115338 161328 115574
rect 161008 115254 161328 115338
rect 161008 115018 161050 115254
rect 161286 115018 161328 115254
rect 161008 114986 161328 115018
rect 114928 111854 115248 111886
rect 114928 111618 114970 111854
rect 115206 111618 115248 111854
rect 114928 111534 115248 111618
rect 114928 111298 114970 111534
rect 115206 111298 115248 111534
rect 114928 111266 115248 111298
rect 145648 111854 145968 111886
rect 145648 111618 145690 111854
rect 145926 111618 145968 111854
rect 145648 111534 145968 111618
rect 145648 111298 145690 111534
rect 145926 111298 145968 111534
rect 145648 111266 145968 111298
rect 176368 111854 176688 111886
rect 176368 111618 176410 111854
rect 176646 111618 176688 111854
rect 176368 111534 176688 111618
rect 176368 111298 176410 111534
rect 176646 111298 176688 111534
rect 176368 111266 176688 111298
rect 189395 98972 189461 98973
rect 189395 98908 189396 98972
rect 189460 98908 189461 98972
rect 189395 98907 189461 98908
rect 96514 97938 96546 98174
rect 96782 97938 96866 98174
rect 97102 97938 97134 98174
rect 96514 97854 97134 97938
rect 96514 97618 96546 97854
rect 96782 97618 96866 97854
rect 97102 97618 97134 97854
rect 92794 58218 92826 58454
rect 93062 58218 93146 58454
rect 93382 58218 93414 58454
rect 92794 58134 93414 58218
rect 92794 57898 92826 58134
rect 93062 57898 93146 58134
rect 93382 57898 93414 58134
rect 92794 22454 93414 57898
rect 92794 22218 92826 22454
rect 93062 22218 93146 22454
rect 93382 22218 93414 22454
rect 92794 22134 93414 22218
rect 92794 21898 92826 22134
rect 93062 21898 93146 22134
rect 93382 21898 93414 22134
rect 89074 -4422 89106 -4186
rect 89342 -4422 89426 -4186
rect 89662 -4422 89694 -4186
rect 89074 -4506 89694 -4422
rect 89074 -4742 89106 -4506
rect 89342 -4742 89426 -4506
rect 89662 -4742 89694 -4506
rect 89074 -7654 89694 -4742
rect 92794 -5146 93414 21898
rect 95006 3773 95066 77742
rect 96514 62174 97134 97618
rect 96514 61938 96546 62174
rect 96782 61938 96866 62174
rect 97102 61938 97134 62174
rect 96514 61854 97134 61938
rect 96514 61618 96546 61854
rect 96782 61618 96866 61854
rect 97102 61618 97134 61854
rect 96514 26174 97134 61618
rect 96514 25938 96546 26174
rect 96782 25938 96866 26174
rect 97102 25938 97134 26174
rect 96514 25854 97134 25938
rect 96514 25618 96546 25854
rect 96782 25618 96866 25854
rect 97102 25618 97134 25854
rect 95003 3772 95069 3773
rect 95003 3708 95004 3772
rect 95068 3708 95069 3772
rect 95003 3707 95069 3708
rect 92794 -5382 92826 -5146
rect 93062 -5382 93146 -5146
rect 93382 -5382 93414 -5146
rect 92794 -5466 93414 -5382
rect 92794 -5702 92826 -5466
rect 93062 -5702 93146 -5466
rect 93382 -5702 93414 -5466
rect 92794 -7654 93414 -5702
rect 96514 -6106 97134 25618
rect 100234 65894 100854 81159
rect 100234 65658 100266 65894
rect 100502 65658 100586 65894
rect 100822 65658 100854 65894
rect 100234 65574 100854 65658
rect 100234 65338 100266 65574
rect 100502 65338 100586 65574
rect 100822 65338 100854 65574
rect 100234 29894 100854 65338
rect 100234 29658 100266 29894
rect 100502 29658 100586 29894
rect 100822 29658 100854 29894
rect 100234 29574 100854 29658
rect 100234 29338 100266 29574
rect 100502 29338 100586 29574
rect 100822 29338 100854 29574
rect 98683 7444 98749 7445
rect 98683 7380 98684 7444
rect 98748 7380 98749 7444
rect 98683 7379 98749 7380
rect 98686 7173 98746 7379
rect 98683 7172 98749 7173
rect 98683 7108 98684 7172
rect 98748 7108 98749 7172
rect 98683 7107 98749 7108
rect 96514 -6342 96546 -6106
rect 96782 -6342 96866 -6106
rect 97102 -6342 97134 -6106
rect 96514 -6426 97134 -6342
rect 96514 -6662 96546 -6426
rect 96782 -6662 96866 -6426
rect 97102 -6662 97134 -6426
rect 96514 -7654 97134 -6662
rect 100234 -7066 100854 29338
rect 100234 -7302 100266 -7066
rect 100502 -7302 100586 -7066
rect 100822 -7302 100854 -7066
rect 100234 -7386 100854 -7302
rect 100234 -7622 100266 -7386
rect 100502 -7622 100586 -7386
rect 100822 -7622 100854 -7386
rect 100234 -7654 100854 -7622
rect 110194 75854 110814 81159
rect 110194 75618 110226 75854
rect 110462 75618 110546 75854
rect 110782 75618 110814 75854
rect 110194 75534 110814 75618
rect 110194 75298 110226 75534
rect 110462 75298 110546 75534
rect 110782 75298 110814 75534
rect 110194 39854 110814 75298
rect 110194 39618 110226 39854
rect 110462 39618 110546 39854
rect 110782 39618 110814 39854
rect 110194 39534 110814 39618
rect 110194 39298 110226 39534
rect 110462 39298 110546 39534
rect 110782 39298 110814 39534
rect 110194 3854 110814 39298
rect 113914 79574 114534 81159
rect 113914 79338 113946 79574
rect 114182 79338 114266 79574
rect 114502 79338 114534 79574
rect 113914 79254 114534 79338
rect 113914 79018 113946 79254
rect 114182 79018 114266 79254
rect 114502 79018 114534 79254
rect 113914 43574 114534 79018
rect 114875 77348 114941 77349
rect 114875 77284 114876 77348
rect 114940 77284 114941 77348
rect 114875 77283 114941 77284
rect 113914 43338 113946 43574
rect 114182 43338 114266 43574
rect 114502 43338 114534 43574
rect 113914 43254 114534 43338
rect 113914 43018 113946 43254
rect 114182 43018 114266 43254
rect 114502 43018 114534 43254
rect 113914 7574 114534 43018
rect 113914 7338 113946 7574
rect 114182 7338 114266 7574
rect 114502 7338 114534 7574
rect 113914 7254 114534 7338
rect 113914 7018 113946 7254
rect 114182 7018 114266 7254
rect 114502 7018 114534 7254
rect 114878 7173 114938 77283
rect 117634 47294 118254 81159
rect 117634 47058 117666 47294
rect 117902 47058 117986 47294
rect 118222 47058 118254 47294
rect 117634 46974 118254 47058
rect 117634 46738 117666 46974
rect 117902 46738 117986 46974
rect 118222 46738 118254 46974
rect 117634 11294 118254 46738
rect 117634 11058 117666 11294
rect 117902 11058 117986 11294
rect 118222 11058 118254 11294
rect 117634 10974 118254 11058
rect 117634 10738 117666 10974
rect 117902 10738 117986 10974
rect 118222 10738 118254 10974
rect 114875 7172 114941 7173
rect 114875 7108 114876 7172
rect 114940 7108 114941 7172
rect 114875 7107 114941 7108
rect 110194 3618 110226 3854
rect 110462 3618 110546 3854
rect 110782 3618 110814 3854
rect 110194 3534 110814 3618
rect 110194 3298 110226 3534
rect 110462 3298 110546 3534
rect 110782 3298 110814 3534
rect 110194 -346 110814 3298
rect 113590 2957 113650 4302
rect 113587 2956 113653 2957
rect 113587 2892 113588 2956
rect 113652 2892 113653 2956
rect 113587 2891 113653 2892
rect 110194 -582 110226 -346
rect 110462 -582 110546 -346
rect 110782 -582 110814 -346
rect 110194 -666 110814 -582
rect 110194 -902 110226 -666
rect 110462 -902 110546 -666
rect 110782 -902 110814 -666
rect 110194 -7654 110814 -902
rect 113914 -1306 114534 7018
rect 113914 -1542 113946 -1306
rect 114182 -1542 114266 -1306
rect 114502 -1542 114534 -1306
rect 113914 -1626 114534 -1542
rect 113914 -1862 113946 -1626
rect 114182 -1862 114266 -1626
rect 114502 -1862 114534 -1626
rect 113914 -7654 114534 -1862
rect 117634 -2266 118254 10738
rect 117634 -2502 117666 -2266
rect 117902 -2502 117986 -2266
rect 118222 -2502 118254 -2266
rect 117634 -2586 118254 -2502
rect 117634 -2822 117666 -2586
rect 117902 -2822 117986 -2586
rect 118222 -2822 118254 -2586
rect 117634 -7654 118254 -2822
rect 121354 51014 121974 81159
rect 121354 50778 121386 51014
rect 121622 50778 121706 51014
rect 121942 50778 121974 51014
rect 121354 50694 121974 50778
rect 121354 50458 121386 50694
rect 121622 50458 121706 50694
rect 121942 50458 121974 50694
rect 121354 15014 121974 50458
rect 121354 14778 121386 15014
rect 121622 14778 121706 15014
rect 121942 14778 121974 15014
rect 121354 14694 121974 14778
rect 121354 14458 121386 14694
rect 121622 14458 121706 14694
rect 121942 14458 121974 14694
rect 121354 -3226 121974 14458
rect 121354 -3462 121386 -3226
rect 121622 -3462 121706 -3226
rect 121942 -3462 121974 -3226
rect 121354 -3546 121974 -3462
rect 121354 -3782 121386 -3546
rect 121622 -3782 121706 -3546
rect 121942 -3782 121974 -3546
rect 121354 -7654 121974 -3782
rect 125074 54734 125694 81159
rect 125074 54498 125106 54734
rect 125342 54498 125426 54734
rect 125662 54498 125694 54734
rect 125074 54414 125694 54498
rect 125074 54178 125106 54414
rect 125342 54178 125426 54414
rect 125662 54178 125694 54414
rect 125074 18734 125694 54178
rect 125074 18498 125106 18734
rect 125342 18498 125426 18734
rect 125662 18498 125694 18734
rect 125074 18414 125694 18498
rect 125074 18178 125106 18414
rect 125342 18178 125426 18414
rect 125662 18178 125694 18414
rect 125074 -4186 125694 18178
rect 125074 -4422 125106 -4186
rect 125342 -4422 125426 -4186
rect 125662 -4422 125694 -4186
rect 125074 -4506 125694 -4422
rect 125074 -4742 125106 -4506
rect 125342 -4742 125426 -4506
rect 125662 -4742 125694 -4506
rect 125074 -7654 125694 -4742
rect 128794 58454 129414 81159
rect 128794 58218 128826 58454
rect 129062 58218 129146 58454
rect 129382 58218 129414 58454
rect 128794 58134 129414 58218
rect 128794 57898 128826 58134
rect 129062 57898 129146 58134
rect 129382 57898 129414 58134
rect 128794 22454 129414 57898
rect 128794 22218 128826 22454
rect 129062 22218 129146 22454
rect 129382 22218 129414 22454
rect 128794 22134 129414 22218
rect 128794 21898 128826 22134
rect 129062 21898 129146 22134
rect 129382 21898 129414 22134
rect 128794 -5146 129414 21898
rect 128794 -5382 128826 -5146
rect 129062 -5382 129146 -5146
rect 129382 -5382 129414 -5146
rect 128794 -5466 129414 -5382
rect 128794 -5702 128826 -5466
rect 129062 -5702 129146 -5466
rect 129382 -5702 129414 -5466
rect 128794 -7654 129414 -5702
rect 132514 62174 133134 81159
rect 132514 61938 132546 62174
rect 132782 61938 132866 62174
rect 133102 61938 133134 62174
rect 132514 61854 133134 61938
rect 132514 61618 132546 61854
rect 132782 61618 132866 61854
rect 133102 61618 133134 61854
rect 132514 26174 133134 61618
rect 132514 25938 132546 26174
rect 132782 25938 132866 26174
rect 133102 25938 133134 26174
rect 132514 25854 133134 25938
rect 132514 25618 132546 25854
rect 132782 25618 132866 25854
rect 133102 25618 133134 25854
rect 132514 -6106 133134 25618
rect 132514 -6342 132546 -6106
rect 132782 -6342 132866 -6106
rect 133102 -6342 133134 -6106
rect 132514 -6426 133134 -6342
rect 132514 -6662 132546 -6426
rect 132782 -6662 132866 -6426
rect 133102 -6662 133134 -6426
rect 132514 -7654 133134 -6662
rect 136234 65894 136854 81159
rect 145051 77892 145117 77893
rect 145051 77828 145052 77892
rect 145116 77828 145117 77892
rect 145051 77827 145117 77828
rect 136234 65658 136266 65894
rect 136502 65658 136586 65894
rect 136822 65658 136854 65894
rect 136234 65574 136854 65658
rect 136234 65338 136266 65574
rect 136502 65338 136586 65574
rect 136822 65338 136854 65574
rect 136234 29894 136854 65338
rect 136234 29658 136266 29894
rect 136502 29658 136586 29894
rect 136822 29658 136854 29894
rect 136234 29574 136854 29658
rect 136234 29338 136266 29574
rect 136502 29338 136586 29574
rect 136822 29338 136854 29574
rect 136234 -7066 136854 29338
rect 145054 9978 145114 77827
rect 146194 75854 146814 81159
rect 146194 75618 146226 75854
rect 146462 75618 146546 75854
rect 146782 75618 146814 75854
rect 146194 75534 146814 75618
rect 146194 75298 146226 75534
rect 146462 75298 146546 75534
rect 146782 75298 146814 75534
rect 146194 39854 146814 75298
rect 146194 39618 146226 39854
rect 146462 39618 146546 39854
rect 146782 39618 146814 39854
rect 146194 39534 146814 39618
rect 146194 39298 146226 39534
rect 146462 39298 146546 39534
rect 146782 39298 146814 39534
rect 136234 -7302 136266 -7066
rect 136502 -7302 136586 -7066
rect 136822 -7302 136854 -7066
rect 136234 -7386 136854 -7302
rect 136234 -7622 136266 -7386
rect 136502 -7622 136586 -7386
rect 136822 -7622 136854 -7386
rect 136234 -7654 136854 -7622
rect 146194 3854 146814 39298
rect 146194 3618 146226 3854
rect 146462 3618 146546 3854
rect 146782 3618 146814 3854
rect 146194 3534 146814 3618
rect 146194 3298 146226 3534
rect 146462 3298 146546 3534
rect 146782 3298 146814 3534
rect 146194 -346 146814 3298
rect 146194 -582 146226 -346
rect 146462 -582 146546 -346
rect 146782 -582 146814 -346
rect 146194 -666 146814 -582
rect 146194 -902 146226 -666
rect 146462 -902 146546 -666
rect 146782 -902 146814 -666
rect 146194 -7654 146814 -902
rect 149914 79574 150534 81159
rect 149914 79338 149946 79574
rect 150182 79338 150266 79574
rect 150502 79338 150534 79574
rect 149914 79254 150534 79338
rect 149914 79018 149946 79254
rect 150182 79018 150266 79254
rect 150502 79018 150534 79254
rect 149914 43574 150534 79018
rect 149914 43338 149946 43574
rect 150182 43338 150266 43574
rect 150502 43338 150534 43574
rect 149914 43254 150534 43338
rect 149914 43018 149946 43254
rect 150182 43018 150266 43254
rect 150502 43018 150534 43254
rect 149914 7574 150534 43018
rect 149914 7338 149946 7574
rect 150182 7338 150266 7574
rect 150502 7338 150534 7574
rect 149914 7254 150534 7338
rect 149914 7018 149946 7254
rect 150182 7018 150266 7254
rect 150502 7018 150534 7254
rect 149914 -1306 150534 7018
rect 149914 -1542 149946 -1306
rect 150182 -1542 150266 -1306
rect 150502 -1542 150534 -1306
rect 149914 -1626 150534 -1542
rect 149914 -1862 149946 -1626
rect 150182 -1862 150266 -1626
rect 150502 -1862 150534 -1626
rect 149914 -7654 150534 -1862
rect 153634 47294 154254 81159
rect 153634 47058 153666 47294
rect 153902 47058 153986 47294
rect 154222 47058 154254 47294
rect 153634 46974 154254 47058
rect 153634 46738 153666 46974
rect 153902 46738 153986 46974
rect 154222 46738 154254 46974
rect 153634 11294 154254 46738
rect 153634 11058 153666 11294
rect 153902 11058 153986 11294
rect 154222 11058 154254 11294
rect 153634 10974 154254 11058
rect 153634 10738 153666 10974
rect 153902 10738 153986 10974
rect 154222 10738 154254 10974
rect 153634 -2266 154254 10738
rect 153634 -2502 153666 -2266
rect 153902 -2502 153986 -2266
rect 154222 -2502 154254 -2266
rect 153634 -2586 154254 -2502
rect 153634 -2822 153666 -2586
rect 153902 -2822 153986 -2586
rect 154222 -2822 154254 -2586
rect 153634 -7654 154254 -2822
rect 157354 51014 157974 81159
rect 157354 50778 157386 51014
rect 157622 50778 157706 51014
rect 157942 50778 157974 51014
rect 157354 50694 157974 50778
rect 157354 50458 157386 50694
rect 157622 50458 157706 50694
rect 157942 50458 157974 50694
rect 157354 15014 157974 50458
rect 157354 14778 157386 15014
rect 157622 14778 157706 15014
rect 157942 14778 157974 15014
rect 157354 14694 157974 14778
rect 157354 14458 157386 14694
rect 157622 14458 157706 14694
rect 157942 14458 157974 14694
rect 157354 -3226 157974 14458
rect 157354 -3462 157386 -3226
rect 157622 -3462 157706 -3226
rect 157942 -3462 157974 -3226
rect 157354 -3546 157974 -3462
rect 157354 -3782 157386 -3546
rect 157622 -3782 157706 -3546
rect 157942 -3782 157974 -3546
rect 157354 -7654 157974 -3782
rect 161074 54734 161694 79988
rect 162899 78164 162965 78165
rect 162899 78100 162900 78164
rect 162964 78100 162965 78164
rect 162899 78099 162965 78100
rect 161074 54498 161106 54734
rect 161342 54498 161426 54734
rect 161662 54498 161694 54734
rect 161074 54414 161694 54498
rect 161074 54178 161106 54414
rect 161342 54178 161426 54414
rect 161662 54178 161694 54414
rect 161074 18734 161694 54178
rect 161074 18498 161106 18734
rect 161342 18498 161426 18734
rect 161662 18498 161694 18734
rect 161074 18414 161694 18498
rect 161074 18178 161106 18414
rect 161342 18178 161426 18414
rect 161662 18178 161694 18414
rect 161074 -4186 161694 18178
rect 162902 8618 162962 78099
rect 164794 58454 165414 81159
rect 164794 58218 164826 58454
rect 165062 58218 165146 58454
rect 165382 58218 165414 58454
rect 164794 58134 165414 58218
rect 164794 57898 164826 58134
rect 165062 57898 165146 58134
rect 165382 57898 165414 58134
rect 164794 22454 165414 57898
rect 164794 22218 164826 22454
rect 165062 22218 165146 22454
rect 165382 22218 165414 22454
rect 164794 22134 165414 22218
rect 164794 21898 164826 22134
rect 165062 21898 165146 22134
rect 165382 21898 165414 22134
rect 161074 -4422 161106 -4186
rect 161342 -4422 161426 -4186
rect 161662 -4422 161694 -4186
rect 161074 -4506 161694 -4422
rect 161074 -4742 161106 -4506
rect 161342 -4742 161426 -4506
rect 161662 -4742 161694 -4506
rect 161074 -7654 161694 -4742
rect 164794 -5146 165414 21898
rect 164794 -5382 164826 -5146
rect 165062 -5382 165146 -5146
rect 165382 -5382 165414 -5146
rect 164794 -5466 165414 -5382
rect 164794 -5702 164826 -5466
rect 165062 -5702 165146 -5466
rect 165382 -5702 165414 -5466
rect 164794 -7654 165414 -5702
rect 168514 62174 169134 81159
rect 168514 61938 168546 62174
rect 168782 61938 168866 62174
rect 169102 61938 169134 62174
rect 168514 61854 169134 61938
rect 168514 61618 168546 61854
rect 168782 61618 168866 61854
rect 169102 61618 169134 61854
rect 168514 26174 169134 61618
rect 168514 25938 168546 26174
rect 168782 25938 168866 26174
rect 169102 25938 169134 26174
rect 168514 25854 169134 25938
rect 168514 25618 168546 25854
rect 168782 25618 168866 25854
rect 169102 25618 169134 25854
rect 168514 -6106 169134 25618
rect 168514 -6342 168546 -6106
rect 168782 -6342 168866 -6106
rect 169102 -6342 169134 -6106
rect 168514 -6426 169134 -6342
rect 168514 -6662 168546 -6426
rect 168782 -6662 168866 -6426
rect 169102 -6662 169134 -6426
rect 168514 -7654 169134 -6662
rect 172234 65894 172854 81159
rect 172234 65658 172266 65894
rect 172502 65658 172586 65894
rect 172822 65658 172854 65894
rect 172234 65574 172854 65658
rect 172234 65338 172266 65574
rect 172502 65338 172586 65574
rect 172822 65338 172854 65574
rect 172234 29894 172854 65338
rect 172234 29658 172266 29894
rect 172502 29658 172586 29894
rect 172822 29658 172854 29894
rect 172234 29574 172854 29658
rect 172234 29338 172266 29574
rect 172502 29338 172586 29574
rect 172822 29338 172854 29574
rect 172234 -7066 172854 29338
rect 173755 7308 173821 7309
rect 173755 7244 173756 7308
rect 173820 7244 173821 7308
rect 173755 7243 173821 7244
rect 173758 6930 173818 7243
rect 173390 6870 173818 6930
rect 173390 3909 173450 6870
rect 177254 4181 177314 77742
rect 182194 75854 182814 81159
rect 182194 75618 182226 75854
rect 182462 75618 182546 75854
rect 182782 75618 182814 75854
rect 182194 75534 182814 75618
rect 182194 75298 182226 75534
rect 182462 75298 182546 75534
rect 182782 75298 182814 75534
rect 182194 39854 182814 75298
rect 182194 39618 182226 39854
rect 182462 39618 182546 39854
rect 182782 39618 182814 39854
rect 182194 39534 182814 39618
rect 182194 39298 182226 39534
rect 182462 39298 182546 39534
rect 182782 39298 182814 39534
rect 177251 4180 177317 4181
rect 177251 4116 177252 4180
rect 177316 4116 177317 4180
rect 177251 4115 177317 4116
rect 173387 3908 173453 3909
rect 173387 3844 173388 3908
rect 173452 3844 173453 3908
rect 173387 3843 173453 3844
rect 182194 3854 182814 39298
rect 172234 -7302 172266 -7066
rect 172502 -7302 172586 -7066
rect 172822 -7302 172854 -7066
rect 172234 -7386 172854 -7302
rect 172234 -7622 172266 -7386
rect 172502 -7622 172586 -7386
rect 172822 -7622 172854 -7386
rect 172234 -7654 172854 -7622
rect 182194 3618 182226 3854
rect 182462 3618 182546 3854
rect 182782 3618 182814 3854
rect 182194 3534 182814 3618
rect 182194 3298 182226 3534
rect 182462 3298 182546 3534
rect 182782 3298 182814 3534
rect 182194 -346 182814 3298
rect 182194 -582 182226 -346
rect 182462 -582 182546 -346
rect 182782 -582 182814 -346
rect 182194 -666 182814 -582
rect 182194 -902 182226 -666
rect 182462 -902 182546 -666
rect 182782 -902 182814 -666
rect 182194 -7654 182814 -902
rect 185914 79574 186534 81159
rect 185914 79338 185946 79574
rect 186182 79338 186266 79574
rect 186502 79338 186534 79574
rect 185914 79254 186534 79338
rect 185914 79018 185946 79254
rect 186182 79018 186266 79254
rect 186502 79018 186534 79254
rect 185914 43574 186534 79018
rect 185914 43338 185946 43574
rect 186182 43338 186266 43574
rect 186502 43338 186534 43574
rect 185914 43254 186534 43338
rect 185914 43018 185946 43254
rect 186182 43018 186266 43254
rect 186502 43018 186534 43254
rect 185914 7574 186534 43018
rect 185914 7338 185946 7574
rect 186182 7338 186266 7574
rect 186502 7338 186534 7574
rect 185914 7254 186534 7338
rect 185914 7018 185946 7254
rect 186182 7018 186266 7254
rect 186502 7018 186534 7254
rect 185914 -1306 186534 7018
rect 189398 4181 189458 98907
rect 189634 83294 190254 118738
rect 190499 114612 190565 114613
rect 190499 114548 190500 114612
rect 190564 114548 190565 114612
rect 190499 114547 190565 114548
rect 189634 83058 189666 83294
rect 189902 83058 189986 83294
rect 190222 83058 190254 83294
rect 189634 82974 190254 83058
rect 189634 82738 189666 82974
rect 189902 82738 189986 82974
rect 190222 82738 190254 82974
rect 189634 47294 190254 82738
rect 189634 47058 189666 47294
rect 189902 47058 189986 47294
rect 190222 47058 190254 47294
rect 189634 46974 190254 47058
rect 189634 46738 189666 46974
rect 189902 46738 189986 46974
rect 190222 46738 190254 46974
rect 189634 11294 190254 46738
rect 190502 16590 190562 114547
rect 190867 92716 190933 92717
rect 190867 92652 190868 92716
rect 190932 92652 190933 92716
rect 190867 92651 190933 92652
rect 190870 16590 190930 92651
rect 191238 16590 191298 127059
rect 190502 16530 190746 16590
rect 190870 16530 191114 16590
rect 191238 16530 191482 16590
rect 189634 11058 189666 11294
rect 189902 11058 189986 11294
rect 190222 11058 190254 11294
rect 189634 10974 190254 11058
rect 189634 10738 189666 10974
rect 189902 10738 189986 10974
rect 190222 10738 190254 10974
rect 189395 4180 189461 4181
rect 189395 4116 189396 4180
rect 189460 4116 189461 4180
rect 189395 4115 189461 4116
rect 185914 -1542 185946 -1306
rect 186182 -1542 186266 -1306
rect 186502 -1542 186534 -1306
rect 185914 -1626 186534 -1542
rect 185914 -1862 185946 -1626
rect 186182 -1862 186266 -1626
rect 186502 -1862 186534 -1626
rect 185914 -7654 186534 -1862
rect 189634 -2266 190254 10738
rect 190686 5898 190746 16530
rect 191054 4045 191114 16530
rect 191422 12018 191482 16530
rect 191790 6930 191850 177107
rect 192342 86461 192402 700435
rect 193354 699014 193974 707162
rect 193354 698778 193386 699014
rect 193622 698778 193706 699014
rect 193942 698778 193974 699014
rect 193354 698694 193974 698778
rect 193354 698458 193386 698694
rect 193622 698458 193706 698694
rect 193942 698458 193974 698694
rect 193354 663014 193974 698458
rect 193354 662778 193386 663014
rect 193622 662778 193706 663014
rect 193942 662778 193974 663014
rect 193354 662694 193974 662778
rect 193354 662458 193386 662694
rect 193622 662458 193706 662694
rect 193942 662458 193974 662694
rect 193354 627014 193974 662458
rect 193354 626778 193386 627014
rect 193622 626778 193706 627014
rect 193942 626778 193974 627014
rect 193354 626694 193974 626778
rect 193354 626458 193386 626694
rect 193622 626458 193706 626694
rect 193942 626458 193974 626694
rect 193354 591014 193974 626458
rect 193354 590778 193386 591014
rect 193622 590778 193706 591014
rect 193942 590778 193974 591014
rect 193354 590694 193974 590778
rect 193354 590458 193386 590694
rect 193622 590458 193706 590694
rect 193942 590458 193974 590694
rect 193354 555014 193974 590458
rect 193354 554778 193386 555014
rect 193622 554778 193706 555014
rect 193942 554778 193974 555014
rect 193354 554694 193974 554778
rect 193354 554458 193386 554694
rect 193622 554458 193706 554694
rect 193942 554458 193974 554694
rect 193354 519014 193974 554458
rect 193354 518778 193386 519014
rect 193622 518778 193706 519014
rect 193942 518778 193974 519014
rect 193354 518694 193974 518778
rect 193354 518458 193386 518694
rect 193622 518458 193706 518694
rect 193942 518458 193974 518694
rect 193354 483014 193974 518458
rect 193354 482778 193386 483014
rect 193622 482778 193706 483014
rect 193942 482778 193974 483014
rect 193354 482694 193974 482778
rect 193354 482458 193386 482694
rect 193622 482458 193706 482694
rect 193942 482458 193974 482694
rect 193354 447014 193974 482458
rect 193354 446778 193386 447014
rect 193622 446778 193706 447014
rect 193942 446778 193974 447014
rect 193354 446694 193974 446778
rect 193354 446458 193386 446694
rect 193622 446458 193706 446694
rect 193942 446458 193974 446694
rect 193354 411014 193974 446458
rect 193354 410778 193386 411014
rect 193622 410778 193706 411014
rect 193942 410778 193974 411014
rect 193354 410694 193974 410778
rect 193354 410458 193386 410694
rect 193622 410458 193706 410694
rect 193942 410458 193974 410694
rect 193354 375014 193974 410458
rect 193354 374778 193386 375014
rect 193622 374778 193706 375014
rect 193942 374778 193974 375014
rect 193354 374694 193974 374778
rect 193354 374458 193386 374694
rect 193622 374458 193706 374694
rect 193942 374458 193974 374694
rect 193354 339014 193974 374458
rect 193354 338778 193386 339014
rect 193622 338778 193706 339014
rect 193942 338778 193974 339014
rect 193354 338694 193974 338778
rect 193354 338458 193386 338694
rect 193622 338458 193706 338694
rect 193942 338458 193974 338694
rect 193354 303014 193974 338458
rect 193354 302778 193386 303014
rect 193622 302778 193706 303014
rect 193942 302778 193974 303014
rect 193354 302694 193974 302778
rect 193354 302458 193386 302694
rect 193622 302458 193706 302694
rect 193942 302458 193974 302694
rect 193354 267014 193974 302458
rect 193354 266778 193386 267014
rect 193622 266778 193706 267014
rect 193942 266778 193974 267014
rect 193354 266694 193974 266778
rect 193354 266458 193386 266694
rect 193622 266458 193706 266694
rect 193942 266458 193974 266694
rect 193354 231014 193974 266458
rect 193354 230778 193386 231014
rect 193622 230778 193706 231014
rect 193942 230778 193974 231014
rect 193354 230694 193974 230778
rect 193354 230458 193386 230694
rect 193622 230458 193706 230694
rect 193942 230458 193974 230694
rect 193354 195014 193974 230458
rect 193354 194778 193386 195014
rect 193622 194778 193706 195014
rect 193942 194778 193974 195014
rect 193354 194694 193974 194778
rect 193354 194458 193386 194694
rect 193622 194458 193706 194694
rect 193942 194458 193974 194694
rect 193354 159014 193974 194458
rect 193354 158778 193386 159014
rect 193622 158778 193706 159014
rect 193942 158778 193974 159014
rect 193354 158694 193974 158778
rect 193354 158458 193386 158694
rect 193622 158458 193706 158694
rect 193942 158458 193974 158694
rect 193354 123014 193974 158458
rect 193354 122778 193386 123014
rect 193622 122778 193706 123014
rect 193942 122778 193974 123014
rect 193354 122694 193974 122778
rect 193354 122458 193386 122694
rect 193622 122458 193706 122694
rect 193942 122458 193974 122694
rect 193354 87014 193974 122458
rect 193354 86778 193386 87014
rect 193622 86778 193706 87014
rect 193942 86778 193974 87014
rect 193354 86694 193974 86778
rect 192339 86460 192405 86461
rect 192339 86396 192340 86460
rect 192404 86396 192405 86460
rect 192339 86395 192405 86396
rect 193354 86458 193386 86694
rect 193622 86458 193706 86694
rect 193942 86458 193974 86694
rect 191971 83332 192037 83333
rect 191971 83268 191972 83332
rect 192036 83268 192037 83332
rect 191971 83267 192037 83268
rect 191974 16590 192034 83267
rect 193354 51014 193974 86458
rect 193354 50778 193386 51014
rect 193622 50778 193706 51014
rect 193942 50778 193974 51014
rect 193354 50694 193974 50778
rect 193354 50458 193386 50694
rect 193622 50458 193706 50694
rect 193942 50458 193974 50694
rect 191974 16530 192218 16590
rect 191422 6870 191850 6930
rect 191422 5218 191482 6870
rect 191790 5813 191850 6342
rect 191787 5812 191853 5813
rect 191787 5748 191788 5812
rect 191852 5748 191853 5812
rect 191787 5747 191853 5748
rect 192158 5541 192218 16530
rect 193354 15014 193974 50458
rect 193354 14778 193386 15014
rect 193622 14778 193706 15014
rect 193942 14778 193974 15014
rect 193354 14694 193974 14778
rect 193354 14458 193386 14694
rect 193622 14458 193706 14694
rect 193942 14458 193974 14694
rect 193075 7444 193141 7445
rect 193075 7380 193076 7444
rect 193140 7380 193141 7444
rect 193075 7379 193141 7380
rect 193078 6901 193138 7379
rect 193075 6900 193141 6901
rect 193075 6836 193076 6900
rect 193140 6836 193141 6900
rect 193075 6835 193141 6836
rect 192155 5540 192221 5541
rect 192155 5476 192156 5540
rect 192220 5476 192221 5540
rect 192155 5475 192221 5476
rect 191051 4044 191117 4045
rect 191051 3980 191052 4044
rect 191116 3980 191117 4044
rect 191051 3979 191117 3980
rect 189634 -2502 189666 -2266
rect 189902 -2502 189986 -2266
rect 190222 -2502 190254 -2266
rect 189634 -2586 190254 -2502
rect 189634 -2822 189666 -2586
rect 189902 -2822 189986 -2586
rect 190222 -2822 190254 -2586
rect 189634 -7654 190254 -2822
rect 193354 -3226 193974 14458
rect 193354 -3462 193386 -3226
rect 193622 -3462 193706 -3226
rect 193942 -3462 193974 -3226
rect 193354 -3546 193974 -3462
rect 193354 -3782 193386 -3546
rect 193622 -3782 193706 -3546
rect 193942 -3782 193974 -3546
rect 193354 -7654 193974 -3782
rect 197074 708678 197694 711590
rect 197074 708442 197106 708678
rect 197342 708442 197426 708678
rect 197662 708442 197694 708678
rect 197074 708358 197694 708442
rect 197074 708122 197106 708358
rect 197342 708122 197426 708358
rect 197662 708122 197694 708358
rect 197074 666734 197694 708122
rect 197074 666498 197106 666734
rect 197342 666498 197426 666734
rect 197662 666498 197694 666734
rect 197074 666414 197694 666498
rect 197074 666178 197106 666414
rect 197342 666178 197426 666414
rect 197662 666178 197694 666414
rect 197074 630734 197694 666178
rect 197074 630498 197106 630734
rect 197342 630498 197426 630734
rect 197662 630498 197694 630734
rect 197074 630414 197694 630498
rect 197074 630178 197106 630414
rect 197342 630178 197426 630414
rect 197662 630178 197694 630414
rect 197074 594734 197694 630178
rect 197074 594498 197106 594734
rect 197342 594498 197426 594734
rect 197662 594498 197694 594734
rect 197074 594414 197694 594498
rect 197074 594178 197106 594414
rect 197342 594178 197426 594414
rect 197662 594178 197694 594414
rect 197074 558734 197694 594178
rect 197074 558498 197106 558734
rect 197342 558498 197426 558734
rect 197662 558498 197694 558734
rect 197074 558414 197694 558498
rect 197074 558178 197106 558414
rect 197342 558178 197426 558414
rect 197662 558178 197694 558414
rect 197074 522734 197694 558178
rect 197074 522498 197106 522734
rect 197342 522498 197426 522734
rect 197662 522498 197694 522734
rect 197074 522414 197694 522498
rect 197074 522178 197106 522414
rect 197342 522178 197426 522414
rect 197662 522178 197694 522414
rect 197074 486734 197694 522178
rect 197074 486498 197106 486734
rect 197342 486498 197426 486734
rect 197662 486498 197694 486734
rect 197074 486414 197694 486498
rect 197074 486178 197106 486414
rect 197342 486178 197426 486414
rect 197662 486178 197694 486414
rect 197074 450734 197694 486178
rect 197074 450498 197106 450734
rect 197342 450498 197426 450734
rect 197662 450498 197694 450734
rect 197074 450414 197694 450498
rect 197074 450178 197106 450414
rect 197342 450178 197426 450414
rect 197662 450178 197694 450414
rect 197074 414734 197694 450178
rect 197074 414498 197106 414734
rect 197342 414498 197426 414734
rect 197662 414498 197694 414734
rect 197074 414414 197694 414498
rect 197074 414178 197106 414414
rect 197342 414178 197426 414414
rect 197662 414178 197694 414414
rect 197074 378734 197694 414178
rect 197074 378498 197106 378734
rect 197342 378498 197426 378734
rect 197662 378498 197694 378734
rect 197074 378414 197694 378498
rect 197074 378178 197106 378414
rect 197342 378178 197426 378414
rect 197662 378178 197694 378414
rect 197074 342734 197694 378178
rect 197074 342498 197106 342734
rect 197342 342498 197426 342734
rect 197662 342498 197694 342734
rect 197074 342414 197694 342498
rect 197074 342178 197106 342414
rect 197342 342178 197426 342414
rect 197662 342178 197694 342414
rect 197074 306734 197694 342178
rect 197074 306498 197106 306734
rect 197342 306498 197426 306734
rect 197662 306498 197694 306734
rect 197074 306414 197694 306498
rect 197074 306178 197106 306414
rect 197342 306178 197426 306414
rect 197662 306178 197694 306414
rect 197074 270734 197694 306178
rect 197074 270498 197106 270734
rect 197342 270498 197426 270734
rect 197662 270498 197694 270734
rect 197074 270414 197694 270498
rect 197074 270178 197106 270414
rect 197342 270178 197426 270414
rect 197662 270178 197694 270414
rect 197074 234734 197694 270178
rect 197074 234498 197106 234734
rect 197342 234498 197426 234734
rect 197662 234498 197694 234734
rect 197074 234414 197694 234498
rect 197074 234178 197106 234414
rect 197342 234178 197426 234414
rect 197662 234178 197694 234414
rect 197074 198734 197694 234178
rect 197074 198498 197106 198734
rect 197342 198498 197426 198734
rect 197662 198498 197694 198734
rect 197074 198414 197694 198498
rect 197074 198178 197106 198414
rect 197342 198178 197426 198414
rect 197662 198178 197694 198414
rect 197074 162734 197694 198178
rect 197074 162498 197106 162734
rect 197342 162498 197426 162734
rect 197662 162498 197694 162734
rect 197074 162414 197694 162498
rect 197074 162178 197106 162414
rect 197342 162178 197426 162414
rect 197662 162178 197694 162414
rect 197074 126734 197694 162178
rect 197074 126498 197106 126734
rect 197342 126498 197426 126734
rect 197662 126498 197694 126734
rect 197074 126414 197694 126498
rect 197074 126178 197106 126414
rect 197342 126178 197426 126414
rect 197662 126178 197694 126414
rect 197074 90734 197694 126178
rect 197074 90498 197106 90734
rect 197342 90498 197426 90734
rect 197662 90498 197694 90734
rect 197074 90414 197694 90498
rect 197074 90178 197106 90414
rect 197342 90178 197426 90414
rect 197662 90178 197694 90414
rect 197074 54734 197694 90178
rect 197074 54498 197106 54734
rect 197342 54498 197426 54734
rect 197662 54498 197694 54734
rect 197074 54414 197694 54498
rect 197074 54178 197106 54414
rect 197342 54178 197426 54414
rect 197662 54178 197694 54414
rect 197074 18734 197694 54178
rect 197074 18498 197106 18734
rect 197342 18498 197426 18734
rect 197662 18498 197694 18734
rect 197074 18414 197694 18498
rect 197074 18178 197106 18414
rect 197342 18178 197426 18414
rect 197662 18178 197694 18414
rect 197074 -4186 197694 18178
rect 197074 -4422 197106 -4186
rect 197342 -4422 197426 -4186
rect 197662 -4422 197694 -4186
rect 197074 -4506 197694 -4422
rect 197074 -4742 197106 -4506
rect 197342 -4742 197426 -4506
rect 197662 -4742 197694 -4506
rect 197074 -7654 197694 -4742
rect 200794 709638 201414 711590
rect 200794 709402 200826 709638
rect 201062 709402 201146 709638
rect 201382 709402 201414 709638
rect 200794 709318 201414 709402
rect 200794 709082 200826 709318
rect 201062 709082 201146 709318
rect 201382 709082 201414 709318
rect 200794 670454 201414 709082
rect 200794 670218 200826 670454
rect 201062 670218 201146 670454
rect 201382 670218 201414 670454
rect 200794 670134 201414 670218
rect 200794 669898 200826 670134
rect 201062 669898 201146 670134
rect 201382 669898 201414 670134
rect 200794 634454 201414 669898
rect 200794 634218 200826 634454
rect 201062 634218 201146 634454
rect 201382 634218 201414 634454
rect 200794 634134 201414 634218
rect 200794 633898 200826 634134
rect 201062 633898 201146 634134
rect 201382 633898 201414 634134
rect 200794 598454 201414 633898
rect 200794 598218 200826 598454
rect 201062 598218 201146 598454
rect 201382 598218 201414 598454
rect 200794 598134 201414 598218
rect 200794 597898 200826 598134
rect 201062 597898 201146 598134
rect 201382 597898 201414 598134
rect 200794 562454 201414 597898
rect 200794 562218 200826 562454
rect 201062 562218 201146 562454
rect 201382 562218 201414 562454
rect 200794 562134 201414 562218
rect 200794 561898 200826 562134
rect 201062 561898 201146 562134
rect 201382 561898 201414 562134
rect 200794 526454 201414 561898
rect 200794 526218 200826 526454
rect 201062 526218 201146 526454
rect 201382 526218 201414 526454
rect 200794 526134 201414 526218
rect 200794 525898 200826 526134
rect 201062 525898 201146 526134
rect 201382 525898 201414 526134
rect 200794 490454 201414 525898
rect 200794 490218 200826 490454
rect 201062 490218 201146 490454
rect 201382 490218 201414 490454
rect 200794 490134 201414 490218
rect 200794 489898 200826 490134
rect 201062 489898 201146 490134
rect 201382 489898 201414 490134
rect 200794 454454 201414 489898
rect 200794 454218 200826 454454
rect 201062 454218 201146 454454
rect 201382 454218 201414 454454
rect 200794 454134 201414 454218
rect 200794 453898 200826 454134
rect 201062 453898 201146 454134
rect 201382 453898 201414 454134
rect 200794 418454 201414 453898
rect 200794 418218 200826 418454
rect 201062 418218 201146 418454
rect 201382 418218 201414 418454
rect 200794 418134 201414 418218
rect 200794 417898 200826 418134
rect 201062 417898 201146 418134
rect 201382 417898 201414 418134
rect 200794 382454 201414 417898
rect 200794 382218 200826 382454
rect 201062 382218 201146 382454
rect 201382 382218 201414 382454
rect 200794 382134 201414 382218
rect 200794 381898 200826 382134
rect 201062 381898 201146 382134
rect 201382 381898 201414 382134
rect 200794 346454 201414 381898
rect 200794 346218 200826 346454
rect 201062 346218 201146 346454
rect 201382 346218 201414 346454
rect 200794 346134 201414 346218
rect 200794 345898 200826 346134
rect 201062 345898 201146 346134
rect 201382 345898 201414 346134
rect 200794 310454 201414 345898
rect 200794 310218 200826 310454
rect 201062 310218 201146 310454
rect 201382 310218 201414 310454
rect 200794 310134 201414 310218
rect 200794 309898 200826 310134
rect 201062 309898 201146 310134
rect 201382 309898 201414 310134
rect 200794 274454 201414 309898
rect 200794 274218 200826 274454
rect 201062 274218 201146 274454
rect 201382 274218 201414 274454
rect 200794 274134 201414 274218
rect 200794 273898 200826 274134
rect 201062 273898 201146 274134
rect 201382 273898 201414 274134
rect 200794 238454 201414 273898
rect 200794 238218 200826 238454
rect 201062 238218 201146 238454
rect 201382 238218 201414 238454
rect 200794 238134 201414 238218
rect 200794 237898 200826 238134
rect 201062 237898 201146 238134
rect 201382 237898 201414 238134
rect 200794 202454 201414 237898
rect 200794 202218 200826 202454
rect 201062 202218 201146 202454
rect 201382 202218 201414 202454
rect 200794 202134 201414 202218
rect 200794 201898 200826 202134
rect 201062 201898 201146 202134
rect 201382 201898 201414 202134
rect 200794 166454 201414 201898
rect 200794 166218 200826 166454
rect 201062 166218 201146 166454
rect 201382 166218 201414 166454
rect 200794 166134 201414 166218
rect 200794 165898 200826 166134
rect 201062 165898 201146 166134
rect 201382 165898 201414 166134
rect 200794 130454 201414 165898
rect 200794 130218 200826 130454
rect 201062 130218 201146 130454
rect 201382 130218 201414 130454
rect 200794 130134 201414 130218
rect 200794 129898 200826 130134
rect 201062 129898 201146 130134
rect 201382 129898 201414 130134
rect 200794 94454 201414 129898
rect 200794 94218 200826 94454
rect 201062 94218 201146 94454
rect 201382 94218 201414 94454
rect 200794 94134 201414 94218
rect 200794 93898 200826 94134
rect 201062 93898 201146 94134
rect 201382 93898 201414 94134
rect 200794 58454 201414 93898
rect 200794 58218 200826 58454
rect 201062 58218 201146 58454
rect 201382 58218 201414 58454
rect 200794 58134 201414 58218
rect 200794 57898 200826 58134
rect 201062 57898 201146 58134
rect 201382 57898 201414 58134
rect 200794 22454 201414 57898
rect 200794 22218 200826 22454
rect 201062 22218 201146 22454
rect 201382 22218 201414 22454
rect 200794 22134 201414 22218
rect 200794 21898 200826 22134
rect 201062 21898 201146 22134
rect 201382 21898 201414 22134
rect 200794 -5146 201414 21898
rect 204514 710598 205134 711590
rect 204514 710362 204546 710598
rect 204782 710362 204866 710598
rect 205102 710362 205134 710598
rect 204514 710278 205134 710362
rect 204514 710042 204546 710278
rect 204782 710042 204866 710278
rect 205102 710042 205134 710278
rect 204514 674174 205134 710042
rect 204514 673938 204546 674174
rect 204782 673938 204866 674174
rect 205102 673938 205134 674174
rect 204514 673854 205134 673938
rect 204514 673618 204546 673854
rect 204782 673618 204866 673854
rect 205102 673618 205134 673854
rect 204514 638174 205134 673618
rect 204514 637938 204546 638174
rect 204782 637938 204866 638174
rect 205102 637938 205134 638174
rect 204514 637854 205134 637938
rect 204514 637618 204546 637854
rect 204782 637618 204866 637854
rect 205102 637618 205134 637854
rect 204514 602174 205134 637618
rect 204514 601938 204546 602174
rect 204782 601938 204866 602174
rect 205102 601938 205134 602174
rect 204514 601854 205134 601938
rect 204514 601618 204546 601854
rect 204782 601618 204866 601854
rect 205102 601618 205134 601854
rect 204514 566174 205134 601618
rect 204514 565938 204546 566174
rect 204782 565938 204866 566174
rect 205102 565938 205134 566174
rect 204514 565854 205134 565938
rect 204514 565618 204546 565854
rect 204782 565618 204866 565854
rect 205102 565618 205134 565854
rect 204514 530174 205134 565618
rect 204514 529938 204546 530174
rect 204782 529938 204866 530174
rect 205102 529938 205134 530174
rect 204514 529854 205134 529938
rect 204514 529618 204546 529854
rect 204782 529618 204866 529854
rect 205102 529618 205134 529854
rect 204514 494174 205134 529618
rect 204514 493938 204546 494174
rect 204782 493938 204866 494174
rect 205102 493938 205134 494174
rect 204514 493854 205134 493938
rect 204514 493618 204546 493854
rect 204782 493618 204866 493854
rect 205102 493618 205134 493854
rect 204514 458174 205134 493618
rect 204514 457938 204546 458174
rect 204782 457938 204866 458174
rect 205102 457938 205134 458174
rect 204514 457854 205134 457938
rect 204514 457618 204546 457854
rect 204782 457618 204866 457854
rect 205102 457618 205134 457854
rect 204514 422174 205134 457618
rect 204514 421938 204546 422174
rect 204782 421938 204866 422174
rect 205102 421938 205134 422174
rect 204514 421854 205134 421938
rect 204514 421618 204546 421854
rect 204782 421618 204866 421854
rect 205102 421618 205134 421854
rect 204514 386174 205134 421618
rect 204514 385938 204546 386174
rect 204782 385938 204866 386174
rect 205102 385938 205134 386174
rect 204514 385854 205134 385938
rect 204514 385618 204546 385854
rect 204782 385618 204866 385854
rect 205102 385618 205134 385854
rect 204514 350174 205134 385618
rect 204514 349938 204546 350174
rect 204782 349938 204866 350174
rect 205102 349938 205134 350174
rect 204514 349854 205134 349938
rect 204514 349618 204546 349854
rect 204782 349618 204866 349854
rect 205102 349618 205134 349854
rect 204514 314174 205134 349618
rect 204514 313938 204546 314174
rect 204782 313938 204866 314174
rect 205102 313938 205134 314174
rect 204514 313854 205134 313938
rect 204514 313618 204546 313854
rect 204782 313618 204866 313854
rect 205102 313618 205134 313854
rect 204514 278174 205134 313618
rect 204514 277938 204546 278174
rect 204782 277938 204866 278174
rect 205102 277938 205134 278174
rect 204514 277854 205134 277938
rect 204514 277618 204546 277854
rect 204782 277618 204866 277854
rect 205102 277618 205134 277854
rect 204514 242174 205134 277618
rect 204514 241938 204546 242174
rect 204782 241938 204866 242174
rect 205102 241938 205134 242174
rect 204514 241854 205134 241938
rect 204514 241618 204546 241854
rect 204782 241618 204866 241854
rect 205102 241618 205134 241854
rect 204514 206174 205134 241618
rect 204514 205938 204546 206174
rect 204782 205938 204866 206174
rect 205102 205938 205134 206174
rect 204514 205854 205134 205938
rect 204514 205618 204546 205854
rect 204782 205618 204866 205854
rect 205102 205618 205134 205854
rect 204514 170174 205134 205618
rect 204514 169938 204546 170174
rect 204782 169938 204866 170174
rect 205102 169938 205134 170174
rect 204514 169854 205134 169938
rect 204514 169618 204546 169854
rect 204782 169618 204866 169854
rect 205102 169618 205134 169854
rect 204514 134174 205134 169618
rect 204514 133938 204546 134174
rect 204782 133938 204866 134174
rect 205102 133938 205134 134174
rect 204514 133854 205134 133938
rect 204514 133618 204546 133854
rect 204782 133618 204866 133854
rect 205102 133618 205134 133854
rect 204514 98174 205134 133618
rect 204514 97938 204546 98174
rect 204782 97938 204866 98174
rect 205102 97938 205134 98174
rect 204514 97854 205134 97938
rect 204514 97618 204546 97854
rect 204782 97618 204866 97854
rect 205102 97618 205134 97854
rect 204514 62174 205134 97618
rect 204514 61938 204546 62174
rect 204782 61938 204866 62174
rect 205102 61938 205134 62174
rect 204514 61854 205134 61938
rect 204514 61618 204546 61854
rect 204782 61618 204866 61854
rect 205102 61618 205134 61854
rect 204514 26174 205134 61618
rect 204514 25938 204546 26174
rect 204782 25938 204866 26174
rect 205102 25938 205134 26174
rect 204514 25854 205134 25938
rect 204514 25618 204546 25854
rect 204782 25618 204866 25854
rect 205102 25618 205134 25854
rect 202827 7444 202893 7445
rect 202827 7380 202828 7444
rect 202892 7380 202893 7444
rect 202827 7379 202893 7380
rect 202830 6930 202890 7379
rect 202646 6901 202890 6930
rect 202643 6900 202890 6901
rect 202643 6836 202644 6900
rect 202708 6870 202890 6900
rect 202708 6836 202709 6870
rect 202643 6835 202709 6836
rect 204118 3229 204178 4302
rect 204115 3228 204181 3229
rect 204115 3164 204116 3228
rect 204180 3164 204181 3228
rect 204115 3163 204181 3164
rect 200794 -5382 200826 -5146
rect 201062 -5382 201146 -5146
rect 201382 -5382 201414 -5146
rect 200794 -5466 201414 -5382
rect 200794 -5702 200826 -5466
rect 201062 -5702 201146 -5466
rect 201382 -5702 201414 -5466
rect 200794 -7654 201414 -5702
rect 204514 -6106 205134 25618
rect 204514 -6342 204546 -6106
rect 204782 -6342 204866 -6106
rect 205102 -6342 205134 -6106
rect 204514 -6426 205134 -6342
rect 204514 -6662 204546 -6426
rect 204782 -6662 204866 -6426
rect 205102 -6662 205134 -6426
rect 204514 -7654 205134 -6662
rect 208234 711558 208854 711590
rect 208234 711322 208266 711558
rect 208502 711322 208586 711558
rect 208822 711322 208854 711558
rect 208234 711238 208854 711322
rect 208234 711002 208266 711238
rect 208502 711002 208586 711238
rect 208822 711002 208854 711238
rect 208234 677894 208854 711002
rect 208234 677658 208266 677894
rect 208502 677658 208586 677894
rect 208822 677658 208854 677894
rect 208234 677574 208854 677658
rect 208234 677338 208266 677574
rect 208502 677338 208586 677574
rect 208822 677338 208854 677574
rect 208234 641894 208854 677338
rect 208234 641658 208266 641894
rect 208502 641658 208586 641894
rect 208822 641658 208854 641894
rect 208234 641574 208854 641658
rect 208234 641338 208266 641574
rect 208502 641338 208586 641574
rect 208822 641338 208854 641574
rect 208234 605894 208854 641338
rect 208234 605658 208266 605894
rect 208502 605658 208586 605894
rect 208822 605658 208854 605894
rect 208234 605574 208854 605658
rect 208234 605338 208266 605574
rect 208502 605338 208586 605574
rect 208822 605338 208854 605574
rect 208234 569894 208854 605338
rect 208234 569658 208266 569894
rect 208502 569658 208586 569894
rect 208822 569658 208854 569894
rect 208234 569574 208854 569658
rect 208234 569338 208266 569574
rect 208502 569338 208586 569574
rect 208822 569338 208854 569574
rect 208234 533894 208854 569338
rect 208234 533658 208266 533894
rect 208502 533658 208586 533894
rect 208822 533658 208854 533894
rect 208234 533574 208854 533658
rect 208234 533338 208266 533574
rect 208502 533338 208586 533574
rect 208822 533338 208854 533574
rect 208234 497894 208854 533338
rect 208234 497658 208266 497894
rect 208502 497658 208586 497894
rect 208822 497658 208854 497894
rect 208234 497574 208854 497658
rect 208234 497338 208266 497574
rect 208502 497338 208586 497574
rect 208822 497338 208854 497574
rect 208234 461894 208854 497338
rect 208234 461658 208266 461894
rect 208502 461658 208586 461894
rect 208822 461658 208854 461894
rect 208234 461574 208854 461658
rect 208234 461338 208266 461574
rect 208502 461338 208586 461574
rect 208822 461338 208854 461574
rect 208234 425894 208854 461338
rect 208234 425658 208266 425894
rect 208502 425658 208586 425894
rect 208822 425658 208854 425894
rect 208234 425574 208854 425658
rect 208234 425338 208266 425574
rect 208502 425338 208586 425574
rect 208822 425338 208854 425574
rect 208234 389894 208854 425338
rect 208234 389658 208266 389894
rect 208502 389658 208586 389894
rect 208822 389658 208854 389894
rect 208234 389574 208854 389658
rect 208234 389338 208266 389574
rect 208502 389338 208586 389574
rect 208822 389338 208854 389574
rect 208234 353894 208854 389338
rect 208234 353658 208266 353894
rect 208502 353658 208586 353894
rect 208822 353658 208854 353894
rect 208234 353574 208854 353658
rect 208234 353338 208266 353574
rect 208502 353338 208586 353574
rect 208822 353338 208854 353574
rect 208234 317894 208854 353338
rect 208234 317658 208266 317894
rect 208502 317658 208586 317894
rect 208822 317658 208854 317894
rect 208234 317574 208854 317658
rect 208234 317338 208266 317574
rect 208502 317338 208586 317574
rect 208822 317338 208854 317574
rect 208234 281894 208854 317338
rect 208234 281658 208266 281894
rect 208502 281658 208586 281894
rect 208822 281658 208854 281894
rect 208234 281574 208854 281658
rect 208234 281338 208266 281574
rect 208502 281338 208586 281574
rect 208822 281338 208854 281574
rect 208234 245894 208854 281338
rect 208234 245658 208266 245894
rect 208502 245658 208586 245894
rect 208822 245658 208854 245894
rect 208234 245574 208854 245658
rect 208234 245338 208266 245574
rect 208502 245338 208586 245574
rect 208822 245338 208854 245574
rect 208234 209894 208854 245338
rect 208234 209658 208266 209894
rect 208502 209658 208586 209894
rect 208822 209658 208854 209894
rect 208234 209574 208854 209658
rect 208234 209338 208266 209574
rect 208502 209338 208586 209574
rect 208822 209338 208854 209574
rect 208234 173894 208854 209338
rect 208234 173658 208266 173894
rect 208502 173658 208586 173894
rect 208822 173658 208854 173894
rect 208234 173574 208854 173658
rect 208234 173338 208266 173574
rect 208502 173338 208586 173574
rect 208822 173338 208854 173574
rect 208234 137894 208854 173338
rect 208234 137658 208266 137894
rect 208502 137658 208586 137894
rect 208822 137658 208854 137894
rect 208234 137574 208854 137658
rect 208234 137338 208266 137574
rect 208502 137338 208586 137574
rect 208822 137338 208854 137574
rect 208234 101894 208854 137338
rect 208234 101658 208266 101894
rect 208502 101658 208586 101894
rect 208822 101658 208854 101894
rect 208234 101574 208854 101658
rect 208234 101338 208266 101574
rect 208502 101338 208586 101574
rect 208822 101338 208854 101574
rect 208234 65894 208854 101338
rect 208234 65658 208266 65894
rect 208502 65658 208586 65894
rect 208822 65658 208854 65894
rect 208234 65574 208854 65658
rect 208234 65338 208266 65574
rect 208502 65338 208586 65574
rect 208822 65338 208854 65574
rect 208234 29894 208854 65338
rect 208234 29658 208266 29894
rect 208502 29658 208586 29894
rect 208822 29658 208854 29894
rect 208234 29574 208854 29658
rect 208234 29338 208266 29574
rect 208502 29338 208586 29574
rect 208822 29338 208854 29574
rect 208234 -7066 208854 29338
rect 218194 704838 218814 711590
rect 218194 704602 218226 704838
rect 218462 704602 218546 704838
rect 218782 704602 218814 704838
rect 218194 704518 218814 704602
rect 218194 704282 218226 704518
rect 218462 704282 218546 704518
rect 218782 704282 218814 704518
rect 218194 687854 218814 704282
rect 218194 687618 218226 687854
rect 218462 687618 218546 687854
rect 218782 687618 218814 687854
rect 218194 687534 218814 687618
rect 218194 687298 218226 687534
rect 218462 687298 218546 687534
rect 218782 687298 218814 687534
rect 218194 651854 218814 687298
rect 218194 651618 218226 651854
rect 218462 651618 218546 651854
rect 218782 651618 218814 651854
rect 218194 651534 218814 651618
rect 218194 651298 218226 651534
rect 218462 651298 218546 651534
rect 218782 651298 218814 651534
rect 218194 615854 218814 651298
rect 218194 615618 218226 615854
rect 218462 615618 218546 615854
rect 218782 615618 218814 615854
rect 218194 615534 218814 615618
rect 218194 615298 218226 615534
rect 218462 615298 218546 615534
rect 218782 615298 218814 615534
rect 218194 579854 218814 615298
rect 218194 579618 218226 579854
rect 218462 579618 218546 579854
rect 218782 579618 218814 579854
rect 218194 579534 218814 579618
rect 218194 579298 218226 579534
rect 218462 579298 218546 579534
rect 218782 579298 218814 579534
rect 218194 543854 218814 579298
rect 218194 543618 218226 543854
rect 218462 543618 218546 543854
rect 218782 543618 218814 543854
rect 218194 543534 218814 543618
rect 218194 543298 218226 543534
rect 218462 543298 218546 543534
rect 218782 543298 218814 543534
rect 218194 507854 218814 543298
rect 218194 507618 218226 507854
rect 218462 507618 218546 507854
rect 218782 507618 218814 507854
rect 218194 507534 218814 507618
rect 218194 507298 218226 507534
rect 218462 507298 218546 507534
rect 218782 507298 218814 507534
rect 218194 471854 218814 507298
rect 218194 471618 218226 471854
rect 218462 471618 218546 471854
rect 218782 471618 218814 471854
rect 218194 471534 218814 471618
rect 218194 471298 218226 471534
rect 218462 471298 218546 471534
rect 218782 471298 218814 471534
rect 218194 435854 218814 471298
rect 218194 435618 218226 435854
rect 218462 435618 218546 435854
rect 218782 435618 218814 435854
rect 218194 435534 218814 435618
rect 218194 435298 218226 435534
rect 218462 435298 218546 435534
rect 218782 435298 218814 435534
rect 218194 399854 218814 435298
rect 218194 399618 218226 399854
rect 218462 399618 218546 399854
rect 218782 399618 218814 399854
rect 218194 399534 218814 399618
rect 218194 399298 218226 399534
rect 218462 399298 218546 399534
rect 218782 399298 218814 399534
rect 218194 363854 218814 399298
rect 218194 363618 218226 363854
rect 218462 363618 218546 363854
rect 218782 363618 218814 363854
rect 218194 363534 218814 363618
rect 218194 363298 218226 363534
rect 218462 363298 218546 363534
rect 218782 363298 218814 363534
rect 218194 327854 218814 363298
rect 218194 327618 218226 327854
rect 218462 327618 218546 327854
rect 218782 327618 218814 327854
rect 218194 327534 218814 327618
rect 218194 327298 218226 327534
rect 218462 327298 218546 327534
rect 218782 327298 218814 327534
rect 218194 291854 218814 327298
rect 218194 291618 218226 291854
rect 218462 291618 218546 291854
rect 218782 291618 218814 291854
rect 218194 291534 218814 291618
rect 218194 291298 218226 291534
rect 218462 291298 218546 291534
rect 218782 291298 218814 291534
rect 218194 255854 218814 291298
rect 218194 255618 218226 255854
rect 218462 255618 218546 255854
rect 218782 255618 218814 255854
rect 218194 255534 218814 255618
rect 218194 255298 218226 255534
rect 218462 255298 218546 255534
rect 218782 255298 218814 255534
rect 218194 219854 218814 255298
rect 218194 219618 218226 219854
rect 218462 219618 218546 219854
rect 218782 219618 218814 219854
rect 218194 219534 218814 219618
rect 218194 219298 218226 219534
rect 218462 219298 218546 219534
rect 218782 219298 218814 219534
rect 218194 183854 218814 219298
rect 218194 183618 218226 183854
rect 218462 183618 218546 183854
rect 218782 183618 218814 183854
rect 218194 183534 218814 183618
rect 218194 183298 218226 183534
rect 218462 183298 218546 183534
rect 218782 183298 218814 183534
rect 218194 147854 218814 183298
rect 218194 147618 218226 147854
rect 218462 147618 218546 147854
rect 218782 147618 218814 147854
rect 218194 147534 218814 147618
rect 218194 147298 218226 147534
rect 218462 147298 218546 147534
rect 218782 147298 218814 147534
rect 218194 111854 218814 147298
rect 218194 111618 218226 111854
rect 218462 111618 218546 111854
rect 218782 111618 218814 111854
rect 218194 111534 218814 111618
rect 218194 111298 218226 111534
rect 218462 111298 218546 111534
rect 218782 111298 218814 111534
rect 218194 75854 218814 111298
rect 218194 75618 218226 75854
rect 218462 75618 218546 75854
rect 218782 75618 218814 75854
rect 218194 75534 218814 75618
rect 218194 75298 218226 75534
rect 218462 75298 218546 75534
rect 218782 75298 218814 75534
rect 218194 39854 218814 75298
rect 218194 39618 218226 39854
rect 218462 39618 218546 39854
rect 218782 39618 218814 39854
rect 218194 39534 218814 39618
rect 218194 39298 218226 39534
rect 218462 39298 218546 39534
rect 218782 39298 218814 39534
rect 212763 7444 212829 7445
rect 212763 7380 212764 7444
rect 212828 7380 212829 7444
rect 212763 7379 212829 7380
rect 212766 6901 212826 7379
rect 212763 6900 212829 6901
rect 212763 6836 212764 6900
rect 212828 6836 212829 6900
rect 212763 6835 212829 6836
rect 208234 -7302 208266 -7066
rect 208502 -7302 208586 -7066
rect 208822 -7302 208854 -7066
rect 208234 -7386 208854 -7302
rect 208234 -7622 208266 -7386
rect 208502 -7622 208586 -7386
rect 208822 -7622 208854 -7386
rect 208234 -7654 208854 -7622
rect 218194 3854 218814 39298
rect 218194 3618 218226 3854
rect 218462 3618 218546 3854
rect 218782 3618 218814 3854
rect 218194 3534 218814 3618
rect 218194 3298 218226 3534
rect 218462 3298 218546 3534
rect 218782 3298 218814 3534
rect 218194 -346 218814 3298
rect 218194 -582 218226 -346
rect 218462 -582 218546 -346
rect 218782 -582 218814 -346
rect 218194 -666 218814 -582
rect 218194 -902 218226 -666
rect 218462 -902 218546 -666
rect 218782 -902 218814 -666
rect 218194 -7654 218814 -902
rect 221914 705798 222534 711590
rect 221914 705562 221946 705798
rect 222182 705562 222266 705798
rect 222502 705562 222534 705798
rect 221914 705478 222534 705562
rect 221914 705242 221946 705478
rect 222182 705242 222266 705478
rect 222502 705242 222534 705478
rect 221914 691574 222534 705242
rect 221914 691338 221946 691574
rect 222182 691338 222266 691574
rect 222502 691338 222534 691574
rect 221914 691254 222534 691338
rect 221914 691018 221946 691254
rect 222182 691018 222266 691254
rect 222502 691018 222534 691254
rect 221914 655574 222534 691018
rect 221914 655338 221946 655574
rect 222182 655338 222266 655574
rect 222502 655338 222534 655574
rect 221914 655254 222534 655338
rect 221914 655018 221946 655254
rect 222182 655018 222266 655254
rect 222502 655018 222534 655254
rect 221914 619574 222534 655018
rect 221914 619338 221946 619574
rect 222182 619338 222266 619574
rect 222502 619338 222534 619574
rect 221914 619254 222534 619338
rect 221914 619018 221946 619254
rect 222182 619018 222266 619254
rect 222502 619018 222534 619254
rect 221914 583574 222534 619018
rect 221914 583338 221946 583574
rect 222182 583338 222266 583574
rect 222502 583338 222534 583574
rect 221914 583254 222534 583338
rect 221914 583018 221946 583254
rect 222182 583018 222266 583254
rect 222502 583018 222534 583254
rect 221914 547574 222534 583018
rect 221914 547338 221946 547574
rect 222182 547338 222266 547574
rect 222502 547338 222534 547574
rect 221914 547254 222534 547338
rect 221914 547018 221946 547254
rect 222182 547018 222266 547254
rect 222502 547018 222534 547254
rect 221914 511574 222534 547018
rect 221914 511338 221946 511574
rect 222182 511338 222266 511574
rect 222502 511338 222534 511574
rect 221914 511254 222534 511338
rect 221914 511018 221946 511254
rect 222182 511018 222266 511254
rect 222502 511018 222534 511254
rect 221914 475574 222534 511018
rect 221914 475338 221946 475574
rect 222182 475338 222266 475574
rect 222502 475338 222534 475574
rect 221914 475254 222534 475338
rect 221914 475018 221946 475254
rect 222182 475018 222266 475254
rect 222502 475018 222534 475254
rect 221914 439574 222534 475018
rect 221914 439338 221946 439574
rect 222182 439338 222266 439574
rect 222502 439338 222534 439574
rect 221914 439254 222534 439338
rect 221914 439018 221946 439254
rect 222182 439018 222266 439254
rect 222502 439018 222534 439254
rect 221914 403574 222534 439018
rect 221914 403338 221946 403574
rect 222182 403338 222266 403574
rect 222502 403338 222534 403574
rect 221914 403254 222534 403338
rect 221914 403018 221946 403254
rect 222182 403018 222266 403254
rect 222502 403018 222534 403254
rect 221914 367574 222534 403018
rect 221914 367338 221946 367574
rect 222182 367338 222266 367574
rect 222502 367338 222534 367574
rect 221914 367254 222534 367338
rect 221914 367018 221946 367254
rect 222182 367018 222266 367254
rect 222502 367018 222534 367254
rect 221914 331574 222534 367018
rect 221914 331338 221946 331574
rect 222182 331338 222266 331574
rect 222502 331338 222534 331574
rect 221914 331254 222534 331338
rect 221914 331018 221946 331254
rect 222182 331018 222266 331254
rect 222502 331018 222534 331254
rect 221914 295574 222534 331018
rect 221914 295338 221946 295574
rect 222182 295338 222266 295574
rect 222502 295338 222534 295574
rect 221914 295254 222534 295338
rect 221914 295018 221946 295254
rect 222182 295018 222266 295254
rect 222502 295018 222534 295254
rect 221914 259574 222534 295018
rect 221914 259338 221946 259574
rect 222182 259338 222266 259574
rect 222502 259338 222534 259574
rect 221914 259254 222534 259338
rect 221914 259018 221946 259254
rect 222182 259018 222266 259254
rect 222502 259018 222534 259254
rect 221914 223574 222534 259018
rect 221914 223338 221946 223574
rect 222182 223338 222266 223574
rect 222502 223338 222534 223574
rect 221914 223254 222534 223338
rect 221914 223018 221946 223254
rect 222182 223018 222266 223254
rect 222502 223018 222534 223254
rect 221914 187574 222534 223018
rect 221914 187338 221946 187574
rect 222182 187338 222266 187574
rect 222502 187338 222534 187574
rect 221914 187254 222534 187338
rect 221914 187018 221946 187254
rect 222182 187018 222266 187254
rect 222502 187018 222534 187254
rect 221914 151574 222534 187018
rect 221914 151338 221946 151574
rect 222182 151338 222266 151574
rect 222502 151338 222534 151574
rect 221914 151254 222534 151338
rect 221914 151018 221946 151254
rect 222182 151018 222266 151254
rect 222502 151018 222534 151254
rect 221914 115574 222534 151018
rect 221914 115338 221946 115574
rect 222182 115338 222266 115574
rect 222502 115338 222534 115574
rect 221914 115254 222534 115338
rect 221914 115018 221946 115254
rect 222182 115018 222266 115254
rect 222502 115018 222534 115254
rect 221914 79574 222534 115018
rect 221914 79338 221946 79574
rect 222182 79338 222266 79574
rect 222502 79338 222534 79574
rect 221914 79254 222534 79338
rect 221914 79018 221946 79254
rect 222182 79018 222266 79254
rect 222502 79018 222534 79254
rect 221914 43574 222534 79018
rect 221914 43338 221946 43574
rect 222182 43338 222266 43574
rect 222502 43338 222534 43574
rect 221914 43254 222534 43338
rect 221914 43018 221946 43254
rect 222182 43018 222266 43254
rect 222502 43018 222534 43254
rect 221914 7574 222534 43018
rect 221914 7338 221946 7574
rect 222182 7338 222266 7574
rect 222502 7338 222534 7574
rect 221914 7254 222534 7338
rect 221914 7018 221946 7254
rect 222182 7018 222266 7254
rect 222502 7018 222534 7254
rect 221914 -1306 222534 7018
rect 221914 -1542 221946 -1306
rect 222182 -1542 222266 -1306
rect 222502 -1542 222534 -1306
rect 221914 -1626 222534 -1542
rect 221914 -1862 221946 -1626
rect 222182 -1862 222266 -1626
rect 222502 -1862 222534 -1626
rect 221914 -7654 222534 -1862
rect 225634 706758 226254 711590
rect 225634 706522 225666 706758
rect 225902 706522 225986 706758
rect 226222 706522 226254 706758
rect 225634 706438 226254 706522
rect 225634 706202 225666 706438
rect 225902 706202 225986 706438
rect 226222 706202 226254 706438
rect 225634 695294 226254 706202
rect 225634 695058 225666 695294
rect 225902 695058 225986 695294
rect 226222 695058 226254 695294
rect 225634 694974 226254 695058
rect 225634 694738 225666 694974
rect 225902 694738 225986 694974
rect 226222 694738 226254 694974
rect 225634 659294 226254 694738
rect 225634 659058 225666 659294
rect 225902 659058 225986 659294
rect 226222 659058 226254 659294
rect 225634 658974 226254 659058
rect 225634 658738 225666 658974
rect 225902 658738 225986 658974
rect 226222 658738 226254 658974
rect 225634 623294 226254 658738
rect 225634 623058 225666 623294
rect 225902 623058 225986 623294
rect 226222 623058 226254 623294
rect 225634 622974 226254 623058
rect 225634 622738 225666 622974
rect 225902 622738 225986 622974
rect 226222 622738 226254 622974
rect 225634 587294 226254 622738
rect 225634 587058 225666 587294
rect 225902 587058 225986 587294
rect 226222 587058 226254 587294
rect 225634 586974 226254 587058
rect 225634 586738 225666 586974
rect 225902 586738 225986 586974
rect 226222 586738 226254 586974
rect 225634 551294 226254 586738
rect 225634 551058 225666 551294
rect 225902 551058 225986 551294
rect 226222 551058 226254 551294
rect 225634 550974 226254 551058
rect 225634 550738 225666 550974
rect 225902 550738 225986 550974
rect 226222 550738 226254 550974
rect 225634 515294 226254 550738
rect 225634 515058 225666 515294
rect 225902 515058 225986 515294
rect 226222 515058 226254 515294
rect 225634 514974 226254 515058
rect 225634 514738 225666 514974
rect 225902 514738 225986 514974
rect 226222 514738 226254 514974
rect 225634 479294 226254 514738
rect 225634 479058 225666 479294
rect 225902 479058 225986 479294
rect 226222 479058 226254 479294
rect 225634 478974 226254 479058
rect 225634 478738 225666 478974
rect 225902 478738 225986 478974
rect 226222 478738 226254 478974
rect 225634 443294 226254 478738
rect 225634 443058 225666 443294
rect 225902 443058 225986 443294
rect 226222 443058 226254 443294
rect 225634 442974 226254 443058
rect 225634 442738 225666 442974
rect 225902 442738 225986 442974
rect 226222 442738 226254 442974
rect 225634 407294 226254 442738
rect 225634 407058 225666 407294
rect 225902 407058 225986 407294
rect 226222 407058 226254 407294
rect 225634 406974 226254 407058
rect 225634 406738 225666 406974
rect 225902 406738 225986 406974
rect 226222 406738 226254 406974
rect 225634 371294 226254 406738
rect 225634 371058 225666 371294
rect 225902 371058 225986 371294
rect 226222 371058 226254 371294
rect 225634 370974 226254 371058
rect 225634 370738 225666 370974
rect 225902 370738 225986 370974
rect 226222 370738 226254 370974
rect 225634 335294 226254 370738
rect 225634 335058 225666 335294
rect 225902 335058 225986 335294
rect 226222 335058 226254 335294
rect 225634 334974 226254 335058
rect 225634 334738 225666 334974
rect 225902 334738 225986 334974
rect 226222 334738 226254 334974
rect 225634 299294 226254 334738
rect 225634 299058 225666 299294
rect 225902 299058 225986 299294
rect 226222 299058 226254 299294
rect 225634 298974 226254 299058
rect 225634 298738 225666 298974
rect 225902 298738 225986 298974
rect 226222 298738 226254 298974
rect 225634 263294 226254 298738
rect 225634 263058 225666 263294
rect 225902 263058 225986 263294
rect 226222 263058 226254 263294
rect 225634 262974 226254 263058
rect 225634 262738 225666 262974
rect 225902 262738 225986 262974
rect 226222 262738 226254 262974
rect 225634 227294 226254 262738
rect 225634 227058 225666 227294
rect 225902 227058 225986 227294
rect 226222 227058 226254 227294
rect 225634 226974 226254 227058
rect 225634 226738 225666 226974
rect 225902 226738 225986 226974
rect 226222 226738 226254 226974
rect 225634 191294 226254 226738
rect 225634 191058 225666 191294
rect 225902 191058 225986 191294
rect 226222 191058 226254 191294
rect 225634 190974 226254 191058
rect 225634 190738 225666 190974
rect 225902 190738 225986 190974
rect 226222 190738 226254 190974
rect 225634 155294 226254 190738
rect 225634 155058 225666 155294
rect 225902 155058 225986 155294
rect 226222 155058 226254 155294
rect 225634 154974 226254 155058
rect 225634 154738 225666 154974
rect 225902 154738 225986 154974
rect 226222 154738 226254 154974
rect 225634 119294 226254 154738
rect 225634 119058 225666 119294
rect 225902 119058 225986 119294
rect 226222 119058 226254 119294
rect 225634 118974 226254 119058
rect 225634 118738 225666 118974
rect 225902 118738 225986 118974
rect 226222 118738 226254 118974
rect 225634 83294 226254 118738
rect 225634 83058 225666 83294
rect 225902 83058 225986 83294
rect 226222 83058 226254 83294
rect 225634 82974 226254 83058
rect 225634 82738 225666 82974
rect 225902 82738 225986 82974
rect 226222 82738 226254 82974
rect 225634 47294 226254 82738
rect 225634 47058 225666 47294
rect 225902 47058 225986 47294
rect 226222 47058 226254 47294
rect 225634 46974 226254 47058
rect 225634 46738 225666 46974
rect 225902 46738 225986 46974
rect 226222 46738 226254 46974
rect 225634 11294 226254 46738
rect 225634 11058 225666 11294
rect 225902 11058 225986 11294
rect 226222 11058 226254 11294
rect 225634 10974 226254 11058
rect 225634 10738 225666 10974
rect 225902 10738 225986 10974
rect 226222 10738 226254 10974
rect 225634 -2266 226254 10738
rect 225634 -2502 225666 -2266
rect 225902 -2502 225986 -2266
rect 226222 -2502 226254 -2266
rect 225634 -2586 226254 -2502
rect 225634 -2822 225666 -2586
rect 225902 -2822 225986 -2586
rect 226222 -2822 226254 -2586
rect 225634 -7654 226254 -2822
rect 229354 707718 229974 711590
rect 229354 707482 229386 707718
rect 229622 707482 229706 707718
rect 229942 707482 229974 707718
rect 229354 707398 229974 707482
rect 229354 707162 229386 707398
rect 229622 707162 229706 707398
rect 229942 707162 229974 707398
rect 229354 699014 229974 707162
rect 229354 698778 229386 699014
rect 229622 698778 229706 699014
rect 229942 698778 229974 699014
rect 229354 698694 229974 698778
rect 229354 698458 229386 698694
rect 229622 698458 229706 698694
rect 229942 698458 229974 698694
rect 229354 663014 229974 698458
rect 229354 662778 229386 663014
rect 229622 662778 229706 663014
rect 229942 662778 229974 663014
rect 229354 662694 229974 662778
rect 229354 662458 229386 662694
rect 229622 662458 229706 662694
rect 229942 662458 229974 662694
rect 229354 627014 229974 662458
rect 229354 626778 229386 627014
rect 229622 626778 229706 627014
rect 229942 626778 229974 627014
rect 229354 626694 229974 626778
rect 229354 626458 229386 626694
rect 229622 626458 229706 626694
rect 229942 626458 229974 626694
rect 229354 591014 229974 626458
rect 229354 590778 229386 591014
rect 229622 590778 229706 591014
rect 229942 590778 229974 591014
rect 229354 590694 229974 590778
rect 229354 590458 229386 590694
rect 229622 590458 229706 590694
rect 229942 590458 229974 590694
rect 229354 555014 229974 590458
rect 229354 554778 229386 555014
rect 229622 554778 229706 555014
rect 229942 554778 229974 555014
rect 229354 554694 229974 554778
rect 229354 554458 229386 554694
rect 229622 554458 229706 554694
rect 229942 554458 229974 554694
rect 229354 519014 229974 554458
rect 229354 518778 229386 519014
rect 229622 518778 229706 519014
rect 229942 518778 229974 519014
rect 229354 518694 229974 518778
rect 229354 518458 229386 518694
rect 229622 518458 229706 518694
rect 229942 518458 229974 518694
rect 229354 483014 229974 518458
rect 229354 482778 229386 483014
rect 229622 482778 229706 483014
rect 229942 482778 229974 483014
rect 229354 482694 229974 482778
rect 229354 482458 229386 482694
rect 229622 482458 229706 482694
rect 229942 482458 229974 482694
rect 229354 447014 229974 482458
rect 229354 446778 229386 447014
rect 229622 446778 229706 447014
rect 229942 446778 229974 447014
rect 229354 446694 229974 446778
rect 229354 446458 229386 446694
rect 229622 446458 229706 446694
rect 229942 446458 229974 446694
rect 229354 411014 229974 446458
rect 229354 410778 229386 411014
rect 229622 410778 229706 411014
rect 229942 410778 229974 411014
rect 229354 410694 229974 410778
rect 229354 410458 229386 410694
rect 229622 410458 229706 410694
rect 229942 410458 229974 410694
rect 229354 375014 229974 410458
rect 229354 374778 229386 375014
rect 229622 374778 229706 375014
rect 229942 374778 229974 375014
rect 229354 374694 229974 374778
rect 229354 374458 229386 374694
rect 229622 374458 229706 374694
rect 229942 374458 229974 374694
rect 229354 339014 229974 374458
rect 229354 338778 229386 339014
rect 229622 338778 229706 339014
rect 229942 338778 229974 339014
rect 229354 338694 229974 338778
rect 229354 338458 229386 338694
rect 229622 338458 229706 338694
rect 229942 338458 229974 338694
rect 229354 303014 229974 338458
rect 229354 302778 229386 303014
rect 229622 302778 229706 303014
rect 229942 302778 229974 303014
rect 229354 302694 229974 302778
rect 229354 302458 229386 302694
rect 229622 302458 229706 302694
rect 229942 302458 229974 302694
rect 229354 267014 229974 302458
rect 229354 266778 229386 267014
rect 229622 266778 229706 267014
rect 229942 266778 229974 267014
rect 229354 266694 229974 266778
rect 229354 266458 229386 266694
rect 229622 266458 229706 266694
rect 229942 266458 229974 266694
rect 229354 231014 229974 266458
rect 229354 230778 229386 231014
rect 229622 230778 229706 231014
rect 229942 230778 229974 231014
rect 229354 230694 229974 230778
rect 229354 230458 229386 230694
rect 229622 230458 229706 230694
rect 229942 230458 229974 230694
rect 229354 195014 229974 230458
rect 229354 194778 229386 195014
rect 229622 194778 229706 195014
rect 229942 194778 229974 195014
rect 229354 194694 229974 194778
rect 229354 194458 229386 194694
rect 229622 194458 229706 194694
rect 229942 194458 229974 194694
rect 229354 159014 229974 194458
rect 229354 158778 229386 159014
rect 229622 158778 229706 159014
rect 229942 158778 229974 159014
rect 229354 158694 229974 158778
rect 229354 158458 229386 158694
rect 229622 158458 229706 158694
rect 229942 158458 229974 158694
rect 229354 123014 229974 158458
rect 229354 122778 229386 123014
rect 229622 122778 229706 123014
rect 229942 122778 229974 123014
rect 229354 122694 229974 122778
rect 229354 122458 229386 122694
rect 229622 122458 229706 122694
rect 229942 122458 229974 122694
rect 229354 87014 229974 122458
rect 229354 86778 229386 87014
rect 229622 86778 229706 87014
rect 229942 86778 229974 87014
rect 229354 86694 229974 86778
rect 229354 86458 229386 86694
rect 229622 86458 229706 86694
rect 229942 86458 229974 86694
rect 229354 51014 229974 86458
rect 229354 50778 229386 51014
rect 229622 50778 229706 51014
rect 229942 50778 229974 51014
rect 229354 50694 229974 50778
rect 229354 50458 229386 50694
rect 229622 50458 229706 50694
rect 229942 50458 229974 50694
rect 229354 15014 229974 50458
rect 229354 14778 229386 15014
rect 229622 14778 229706 15014
rect 229942 14778 229974 15014
rect 229354 14694 229974 14778
rect 229354 14458 229386 14694
rect 229622 14458 229706 14694
rect 229942 14458 229974 14694
rect 229354 -3226 229974 14458
rect 229354 -3462 229386 -3226
rect 229622 -3462 229706 -3226
rect 229942 -3462 229974 -3226
rect 229354 -3546 229974 -3462
rect 229354 -3782 229386 -3546
rect 229622 -3782 229706 -3546
rect 229942 -3782 229974 -3546
rect 229354 -7654 229974 -3782
rect 233074 708678 233694 711590
rect 233074 708442 233106 708678
rect 233342 708442 233426 708678
rect 233662 708442 233694 708678
rect 233074 708358 233694 708442
rect 233074 708122 233106 708358
rect 233342 708122 233426 708358
rect 233662 708122 233694 708358
rect 233074 666734 233694 708122
rect 233074 666498 233106 666734
rect 233342 666498 233426 666734
rect 233662 666498 233694 666734
rect 233074 666414 233694 666498
rect 233074 666178 233106 666414
rect 233342 666178 233426 666414
rect 233662 666178 233694 666414
rect 233074 630734 233694 666178
rect 233074 630498 233106 630734
rect 233342 630498 233426 630734
rect 233662 630498 233694 630734
rect 233074 630414 233694 630498
rect 233074 630178 233106 630414
rect 233342 630178 233426 630414
rect 233662 630178 233694 630414
rect 233074 594734 233694 630178
rect 233074 594498 233106 594734
rect 233342 594498 233426 594734
rect 233662 594498 233694 594734
rect 233074 594414 233694 594498
rect 233074 594178 233106 594414
rect 233342 594178 233426 594414
rect 233662 594178 233694 594414
rect 233074 558734 233694 594178
rect 233074 558498 233106 558734
rect 233342 558498 233426 558734
rect 233662 558498 233694 558734
rect 233074 558414 233694 558498
rect 233074 558178 233106 558414
rect 233342 558178 233426 558414
rect 233662 558178 233694 558414
rect 233074 522734 233694 558178
rect 233074 522498 233106 522734
rect 233342 522498 233426 522734
rect 233662 522498 233694 522734
rect 233074 522414 233694 522498
rect 233074 522178 233106 522414
rect 233342 522178 233426 522414
rect 233662 522178 233694 522414
rect 233074 486734 233694 522178
rect 233074 486498 233106 486734
rect 233342 486498 233426 486734
rect 233662 486498 233694 486734
rect 233074 486414 233694 486498
rect 233074 486178 233106 486414
rect 233342 486178 233426 486414
rect 233662 486178 233694 486414
rect 233074 450734 233694 486178
rect 233074 450498 233106 450734
rect 233342 450498 233426 450734
rect 233662 450498 233694 450734
rect 233074 450414 233694 450498
rect 233074 450178 233106 450414
rect 233342 450178 233426 450414
rect 233662 450178 233694 450414
rect 233074 414734 233694 450178
rect 233074 414498 233106 414734
rect 233342 414498 233426 414734
rect 233662 414498 233694 414734
rect 233074 414414 233694 414498
rect 233074 414178 233106 414414
rect 233342 414178 233426 414414
rect 233662 414178 233694 414414
rect 233074 378734 233694 414178
rect 233074 378498 233106 378734
rect 233342 378498 233426 378734
rect 233662 378498 233694 378734
rect 233074 378414 233694 378498
rect 233074 378178 233106 378414
rect 233342 378178 233426 378414
rect 233662 378178 233694 378414
rect 233074 342734 233694 378178
rect 233074 342498 233106 342734
rect 233342 342498 233426 342734
rect 233662 342498 233694 342734
rect 233074 342414 233694 342498
rect 233074 342178 233106 342414
rect 233342 342178 233426 342414
rect 233662 342178 233694 342414
rect 233074 306734 233694 342178
rect 233074 306498 233106 306734
rect 233342 306498 233426 306734
rect 233662 306498 233694 306734
rect 233074 306414 233694 306498
rect 233074 306178 233106 306414
rect 233342 306178 233426 306414
rect 233662 306178 233694 306414
rect 233074 270734 233694 306178
rect 233074 270498 233106 270734
rect 233342 270498 233426 270734
rect 233662 270498 233694 270734
rect 233074 270414 233694 270498
rect 233074 270178 233106 270414
rect 233342 270178 233426 270414
rect 233662 270178 233694 270414
rect 233074 234734 233694 270178
rect 233074 234498 233106 234734
rect 233342 234498 233426 234734
rect 233662 234498 233694 234734
rect 233074 234414 233694 234498
rect 233074 234178 233106 234414
rect 233342 234178 233426 234414
rect 233662 234178 233694 234414
rect 233074 198734 233694 234178
rect 233074 198498 233106 198734
rect 233342 198498 233426 198734
rect 233662 198498 233694 198734
rect 233074 198414 233694 198498
rect 233074 198178 233106 198414
rect 233342 198178 233426 198414
rect 233662 198178 233694 198414
rect 233074 162734 233694 198178
rect 233074 162498 233106 162734
rect 233342 162498 233426 162734
rect 233662 162498 233694 162734
rect 233074 162414 233694 162498
rect 233074 162178 233106 162414
rect 233342 162178 233426 162414
rect 233662 162178 233694 162414
rect 233074 126734 233694 162178
rect 233074 126498 233106 126734
rect 233342 126498 233426 126734
rect 233662 126498 233694 126734
rect 233074 126414 233694 126498
rect 233074 126178 233106 126414
rect 233342 126178 233426 126414
rect 233662 126178 233694 126414
rect 233074 90734 233694 126178
rect 233074 90498 233106 90734
rect 233342 90498 233426 90734
rect 233662 90498 233694 90734
rect 233074 90414 233694 90498
rect 233074 90178 233106 90414
rect 233342 90178 233426 90414
rect 233662 90178 233694 90414
rect 233074 54734 233694 90178
rect 233074 54498 233106 54734
rect 233342 54498 233426 54734
rect 233662 54498 233694 54734
rect 233074 54414 233694 54498
rect 233074 54178 233106 54414
rect 233342 54178 233426 54414
rect 233662 54178 233694 54414
rect 233074 18734 233694 54178
rect 233074 18498 233106 18734
rect 233342 18498 233426 18734
rect 233662 18498 233694 18734
rect 233074 18414 233694 18498
rect 233074 18178 233106 18414
rect 233342 18178 233426 18414
rect 233662 18178 233694 18414
rect 233074 -4186 233694 18178
rect 233074 -4422 233106 -4186
rect 233342 -4422 233426 -4186
rect 233662 -4422 233694 -4186
rect 233074 -4506 233694 -4422
rect 233074 -4742 233106 -4506
rect 233342 -4742 233426 -4506
rect 233662 -4742 233694 -4506
rect 233074 -7654 233694 -4742
rect 236794 709638 237414 711590
rect 236794 709402 236826 709638
rect 237062 709402 237146 709638
rect 237382 709402 237414 709638
rect 236794 709318 237414 709402
rect 236794 709082 236826 709318
rect 237062 709082 237146 709318
rect 237382 709082 237414 709318
rect 236794 670454 237414 709082
rect 236794 670218 236826 670454
rect 237062 670218 237146 670454
rect 237382 670218 237414 670454
rect 236794 670134 237414 670218
rect 236794 669898 236826 670134
rect 237062 669898 237146 670134
rect 237382 669898 237414 670134
rect 236794 634454 237414 669898
rect 236794 634218 236826 634454
rect 237062 634218 237146 634454
rect 237382 634218 237414 634454
rect 236794 634134 237414 634218
rect 236794 633898 236826 634134
rect 237062 633898 237146 634134
rect 237382 633898 237414 634134
rect 236794 598454 237414 633898
rect 236794 598218 236826 598454
rect 237062 598218 237146 598454
rect 237382 598218 237414 598454
rect 236794 598134 237414 598218
rect 236794 597898 236826 598134
rect 237062 597898 237146 598134
rect 237382 597898 237414 598134
rect 236794 562454 237414 597898
rect 236794 562218 236826 562454
rect 237062 562218 237146 562454
rect 237382 562218 237414 562454
rect 236794 562134 237414 562218
rect 236794 561898 236826 562134
rect 237062 561898 237146 562134
rect 237382 561898 237414 562134
rect 236794 526454 237414 561898
rect 236794 526218 236826 526454
rect 237062 526218 237146 526454
rect 237382 526218 237414 526454
rect 236794 526134 237414 526218
rect 236794 525898 236826 526134
rect 237062 525898 237146 526134
rect 237382 525898 237414 526134
rect 236794 490454 237414 525898
rect 236794 490218 236826 490454
rect 237062 490218 237146 490454
rect 237382 490218 237414 490454
rect 236794 490134 237414 490218
rect 236794 489898 236826 490134
rect 237062 489898 237146 490134
rect 237382 489898 237414 490134
rect 236794 454454 237414 489898
rect 236794 454218 236826 454454
rect 237062 454218 237146 454454
rect 237382 454218 237414 454454
rect 236794 454134 237414 454218
rect 236794 453898 236826 454134
rect 237062 453898 237146 454134
rect 237382 453898 237414 454134
rect 236794 418454 237414 453898
rect 236794 418218 236826 418454
rect 237062 418218 237146 418454
rect 237382 418218 237414 418454
rect 236794 418134 237414 418218
rect 236794 417898 236826 418134
rect 237062 417898 237146 418134
rect 237382 417898 237414 418134
rect 236794 382454 237414 417898
rect 236794 382218 236826 382454
rect 237062 382218 237146 382454
rect 237382 382218 237414 382454
rect 236794 382134 237414 382218
rect 236794 381898 236826 382134
rect 237062 381898 237146 382134
rect 237382 381898 237414 382134
rect 236794 346454 237414 381898
rect 236794 346218 236826 346454
rect 237062 346218 237146 346454
rect 237382 346218 237414 346454
rect 236794 346134 237414 346218
rect 236794 345898 236826 346134
rect 237062 345898 237146 346134
rect 237382 345898 237414 346134
rect 236794 310454 237414 345898
rect 236794 310218 236826 310454
rect 237062 310218 237146 310454
rect 237382 310218 237414 310454
rect 236794 310134 237414 310218
rect 236794 309898 236826 310134
rect 237062 309898 237146 310134
rect 237382 309898 237414 310134
rect 236794 274454 237414 309898
rect 236794 274218 236826 274454
rect 237062 274218 237146 274454
rect 237382 274218 237414 274454
rect 236794 274134 237414 274218
rect 236794 273898 236826 274134
rect 237062 273898 237146 274134
rect 237382 273898 237414 274134
rect 236794 238454 237414 273898
rect 236794 238218 236826 238454
rect 237062 238218 237146 238454
rect 237382 238218 237414 238454
rect 236794 238134 237414 238218
rect 236794 237898 236826 238134
rect 237062 237898 237146 238134
rect 237382 237898 237414 238134
rect 236794 202454 237414 237898
rect 236794 202218 236826 202454
rect 237062 202218 237146 202454
rect 237382 202218 237414 202454
rect 236794 202134 237414 202218
rect 236794 201898 236826 202134
rect 237062 201898 237146 202134
rect 237382 201898 237414 202134
rect 236794 166454 237414 201898
rect 236794 166218 236826 166454
rect 237062 166218 237146 166454
rect 237382 166218 237414 166454
rect 236794 166134 237414 166218
rect 236794 165898 236826 166134
rect 237062 165898 237146 166134
rect 237382 165898 237414 166134
rect 236794 130454 237414 165898
rect 236794 130218 236826 130454
rect 237062 130218 237146 130454
rect 237382 130218 237414 130454
rect 236794 130134 237414 130218
rect 236794 129898 236826 130134
rect 237062 129898 237146 130134
rect 237382 129898 237414 130134
rect 236794 94454 237414 129898
rect 236794 94218 236826 94454
rect 237062 94218 237146 94454
rect 237382 94218 237414 94454
rect 236794 94134 237414 94218
rect 236794 93898 236826 94134
rect 237062 93898 237146 94134
rect 237382 93898 237414 94134
rect 236794 58454 237414 93898
rect 236794 58218 236826 58454
rect 237062 58218 237146 58454
rect 237382 58218 237414 58454
rect 236794 58134 237414 58218
rect 236794 57898 236826 58134
rect 237062 57898 237146 58134
rect 237382 57898 237414 58134
rect 236794 22454 237414 57898
rect 236794 22218 236826 22454
rect 237062 22218 237146 22454
rect 237382 22218 237414 22454
rect 236794 22134 237414 22218
rect 236794 21898 236826 22134
rect 237062 21898 237146 22134
rect 237382 21898 237414 22134
rect 236794 -5146 237414 21898
rect 236794 -5382 236826 -5146
rect 237062 -5382 237146 -5146
rect 237382 -5382 237414 -5146
rect 236794 -5466 237414 -5382
rect 236794 -5702 236826 -5466
rect 237062 -5702 237146 -5466
rect 237382 -5702 237414 -5466
rect 236794 -7654 237414 -5702
rect 240514 710598 241134 711590
rect 240514 710362 240546 710598
rect 240782 710362 240866 710598
rect 241102 710362 241134 710598
rect 240514 710278 241134 710362
rect 240514 710042 240546 710278
rect 240782 710042 240866 710278
rect 241102 710042 241134 710278
rect 240514 674174 241134 710042
rect 240514 673938 240546 674174
rect 240782 673938 240866 674174
rect 241102 673938 241134 674174
rect 240514 673854 241134 673938
rect 240514 673618 240546 673854
rect 240782 673618 240866 673854
rect 241102 673618 241134 673854
rect 240514 638174 241134 673618
rect 240514 637938 240546 638174
rect 240782 637938 240866 638174
rect 241102 637938 241134 638174
rect 240514 637854 241134 637938
rect 240514 637618 240546 637854
rect 240782 637618 240866 637854
rect 241102 637618 241134 637854
rect 240514 602174 241134 637618
rect 240514 601938 240546 602174
rect 240782 601938 240866 602174
rect 241102 601938 241134 602174
rect 240514 601854 241134 601938
rect 240514 601618 240546 601854
rect 240782 601618 240866 601854
rect 241102 601618 241134 601854
rect 240514 566174 241134 601618
rect 240514 565938 240546 566174
rect 240782 565938 240866 566174
rect 241102 565938 241134 566174
rect 240514 565854 241134 565938
rect 240514 565618 240546 565854
rect 240782 565618 240866 565854
rect 241102 565618 241134 565854
rect 240514 530174 241134 565618
rect 240514 529938 240546 530174
rect 240782 529938 240866 530174
rect 241102 529938 241134 530174
rect 240514 529854 241134 529938
rect 240514 529618 240546 529854
rect 240782 529618 240866 529854
rect 241102 529618 241134 529854
rect 240514 494174 241134 529618
rect 240514 493938 240546 494174
rect 240782 493938 240866 494174
rect 241102 493938 241134 494174
rect 240514 493854 241134 493938
rect 240514 493618 240546 493854
rect 240782 493618 240866 493854
rect 241102 493618 241134 493854
rect 240514 458174 241134 493618
rect 240514 457938 240546 458174
rect 240782 457938 240866 458174
rect 241102 457938 241134 458174
rect 240514 457854 241134 457938
rect 240514 457618 240546 457854
rect 240782 457618 240866 457854
rect 241102 457618 241134 457854
rect 240514 422174 241134 457618
rect 240514 421938 240546 422174
rect 240782 421938 240866 422174
rect 241102 421938 241134 422174
rect 240514 421854 241134 421938
rect 240514 421618 240546 421854
rect 240782 421618 240866 421854
rect 241102 421618 241134 421854
rect 240514 386174 241134 421618
rect 240514 385938 240546 386174
rect 240782 385938 240866 386174
rect 241102 385938 241134 386174
rect 240514 385854 241134 385938
rect 240514 385618 240546 385854
rect 240782 385618 240866 385854
rect 241102 385618 241134 385854
rect 240514 350174 241134 385618
rect 240514 349938 240546 350174
rect 240782 349938 240866 350174
rect 241102 349938 241134 350174
rect 240514 349854 241134 349938
rect 240514 349618 240546 349854
rect 240782 349618 240866 349854
rect 241102 349618 241134 349854
rect 240514 314174 241134 349618
rect 240514 313938 240546 314174
rect 240782 313938 240866 314174
rect 241102 313938 241134 314174
rect 240514 313854 241134 313938
rect 240514 313618 240546 313854
rect 240782 313618 240866 313854
rect 241102 313618 241134 313854
rect 240514 278174 241134 313618
rect 240514 277938 240546 278174
rect 240782 277938 240866 278174
rect 241102 277938 241134 278174
rect 240514 277854 241134 277938
rect 240514 277618 240546 277854
rect 240782 277618 240866 277854
rect 241102 277618 241134 277854
rect 240514 242174 241134 277618
rect 240514 241938 240546 242174
rect 240782 241938 240866 242174
rect 241102 241938 241134 242174
rect 240514 241854 241134 241938
rect 240514 241618 240546 241854
rect 240782 241618 240866 241854
rect 241102 241618 241134 241854
rect 240514 206174 241134 241618
rect 240514 205938 240546 206174
rect 240782 205938 240866 206174
rect 241102 205938 241134 206174
rect 240514 205854 241134 205938
rect 240514 205618 240546 205854
rect 240782 205618 240866 205854
rect 241102 205618 241134 205854
rect 240514 170174 241134 205618
rect 240514 169938 240546 170174
rect 240782 169938 240866 170174
rect 241102 169938 241134 170174
rect 240514 169854 241134 169938
rect 240514 169618 240546 169854
rect 240782 169618 240866 169854
rect 241102 169618 241134 169854
rect 240514 134174 241134 169618
rect 240514 133938 240546 134174
rect 240782 133938 240866 134174
rect 241102 133938 241134 134174
rect 240514 133854 241134 133938
rect 240514 133618 240546 133854
rect 240782 133618 240866 133854
rect 241102 133618 241134 133854
rect 240514 98174 241134 133618
rect 240514 97938 240546 98174
rect 240782 97938 240866 98174
rect 241102 97938 241134 98174
rect 240514 97854 241134 97938
rect 240514 97618 240546 97854
rect 240782 97618 240866 97854
rect 241102 97618 241134 97854
rect 240514 62174 241134 97618
rect 240514 61938 240546 62174
rect 240782 61938 240866 62174
rect 241102 61938 241134 62174
rect 240514 61854 241134 61938
rect 240514 61618 240546 61854
rect 240782 61618 240866 61854
rect 241102 61618 241134 61854
rect 240514 26174 241134 61618
rect 240514 25938 240546 26174
rect 240782 25938 240866 26174
rect 241102 25938 241134 26174
rect 240514 25854 241134 25938
rect 240514 25618 240546 25854
rect 240782 25618 240866 25854
rect 241102 25618 241134 25854
rect 240514 -6106 241134 25618
rect 244234 711558 244854 711590
rect 244234 711322 244266 711558
rect 244502 711322 244586 711558
rect 244822 711322 244854 711558
rect 244234 711238 244854 711322
rect 244234 711002 244266 711238
rect 244502 711002 244586 711238
rect 244822 711002 244854 711238
rect 244234 677894 244854 711002
rect 244234 677658 244266 677894
rect 244502 677658 244586 677894
rect 244822 677658 244854 677894
rect 244234 677574 244854 677658
rect 244234 677338 244266 677574
rect 244502 677338 244586 677574
rect 244822 677338 244854 677574
rect 244234 641894 244854 677338
rect 244234 641658 244266 641894
rect 244502 641658 244586 641894
rect 244822 641658 244854 641894
rect 244234 641574 244854 641658
rect 244234 641338 244266 641574
rect 244502 641338 244586 641574
rect 244822 641338 244854 641574
rect 244234 605894 244854 641338
rect 244234 605658 244266 605894
rect 244502 605658 244586 605894
rect 244822 605658 244854 605894
rect 244234 605574 244854 605658
rect 244234 605338 244266 605574
rect 244502 605338 244586 605574
rect 244822 605338 244854 605574
rect 244234 569894 244854 605338
rect 244234 569658 244266 569894
rect 244502 569658 244586 569894
rect 244822 569658 244854 569894
rect 244234 569574 244854 569658
rect 244234 569338 244266 569574
rect 244502 569338 244586 569574
rect 244822 569338 244854 569574
rect 244234 533894 244854 569338
rect 244234 533658 244266 533894
rect 244502 533658 244586 533894
rect 244822 533658 244854 533894
rect 244234 533574 244854 533658
rect 244234 533338 244266 533574
rect 244502 533338 244586 533574
rect 244822 533338 244854 533574
rect 244234 497894 244854 533338
rect 244234 497658 244266 497894
rect 244502 497658 244586 497894
rect 244822 497658 244854 497894
rect 244234 497574 244854 497658
rect 244234 497338 244266 497574
rect 244502 497338 244586 497574
rect 244822 497338 244854 497574
rect 244234 461894 244854 497338
rect 244234 461658 244266 461894
rect 244502 461658 244586 461894
rect 244822 461658 244854 461894
rect 244234 461574 244854 461658
rect 244234 461338 244266 461574
rect 244502 461338 244586 461574
rect 244822 461338 244854 461574
rect 244234 425894 244854 461338
rect 244234 425658 244266 425894
rect 244502 425658 244586 425894
rect 244822 425658 244854 425894
rect 244234 425574 244854 425658
rect 244234 425338 244266 425574
rect 244502 425338 244586 425574
rect 244822 425338 244854 425574
rect 244234 389894 244854 425338
rect 244234 389658 244266 389894
rect 244502 389658 244586 389894
rect 244822 389658 244854 389894
rect 244234 389574 244854 389658
rect 244234 389338 244266 389574
rect 244502 389338 244586 389574
rect 244822 389338 244854 389574
rect 244234 353894 244854 389338
rect 244234 353658 244266 353894
rect 244502 353658 244586 353894
rect 244822 353658 244854 353894
rect 244234 353574 244854 353658
rect 244234 353338 244266 353574
rect 244502 353338 244586 353574
rect 244822 353338 244854 353574
rect 244234 317894 244854 353338
rect 244234 317658 244266 317894
rect 244502 317658 244586 317894
rect 244822 317658 244854 317894
rect 244234 317574 244854 317658
rect 244234 317338 244266 317574
rect 244502 317338 244586 317574
rect 244822 317338 244854 317574
rect 244234 281894 244854 317338
rect 244234 281658 244266 281894
rect 244502 281658 244586 281894
rect 244822 281658 244854 281894
rect 244234 281574 244854 281658
rect 244234 281338 244266 281574
rect 244502 281338 244586 281574
rect 244822 281338 244854 281574
rect 244234 245894 244854 281338
rect 244234 245658 244266 245894
rect 244502 245658 244586 245894
rect 244822 245658 244854 245894
rect 244234 245574 244854 245658
rect 244234 245338 244266 245574
rect 244502 245338 244586 245574
rect 244822 245338 244854 245574
rect 244234 209894 244854 245338
rect 244234 209658 244266 209894
rect 244502 209658 244586 209894
rect 244822 209658 244854 209894
rect 244234 209574 244854 209658
rect 244234 209338 244266 209574
rect 244502 209338 244586 209574
rect 244822 209338 244854 209574
rect 244234 173894 244854 209338
rect 244234 173658 244266 173894
rect 244502 173658 244586 173894
rect 244822 173658 244854 173894
rect 244234 173574 244854 173658
rect 244234 173338 244266 173574
rect 244502 173338 244586 173574
rect 244822 173338 244854 173574
rect 244234 137894 244854 173338
rect 244234 137658 244266 137894
rect 244502 137658 244586 137894
rect 244822 137658 244854 137894
rect 244234 137574 244854 137658
rect 244234 137338 244266 137574
rect 244502 137338 244586 137574
rect 244822 137338 244854 137574
rect 244234 101894 244854 137338
rect 244234 101658 244266 101894
rect 244502 101658 244586 101894
rect 244822 101658 244854 101894
rect 244234 101574 244854 101658
rect 244234 101338 244266 101574
rect 244502 101338 244586 101574
rect 244822 101338 244854 101574
rect 244234 65894 244854 101338
rect 244234 65658 244266 65894
rect 244502 65658 244586 65894
rect 244822 65658 244854 65894
rect 244234 65574 244854 65658
rect 244234 65338 244266 65574
rect 244502 65338 244586 65574
rect 244822 65338 244854 65574
rect 244234 29894 244854 65338
rect 244234 29658 244266 29894
rect 244502 29658 244586 29894
rect 244822 29658 244854 29894
rect 244234 29574 244854 29658
rect 244234 29338 244266 29574
rect 244502 29338 244586 29574
rect 244822 29338 244854 29574
rect 243491 7444 243557 7445
rect 243491 7380 243492 7444
rect 243556 7380 243557 7444
rect 243491 7379 243557 7380
rect 243494 7173 243554 7379
rect 243491 7172 243557 7173
rect 243491 7108 243492 7172
rect 243556 7108 243557 7172
rect 243491 7107 243557 7108
rect 240514 -6342 240546 -6106
rect 240782 -6342 240866 -6106
rect 241102 -6342 241134 -6106
rect 240514 -6426 241134 -6342
rect 240514 -6662 240546 -6426
rect 240782 -6662 240866 -6426
rect 241102 -6662 241134 -6426
rect 240514 -7654 241134 -6662
rect 244234 -7066 244854 29338
rect 244234 -7302 244266 -7066
rect 244502 -7302 244586 -7066
rect 244822 -7302 244854 -7066
rect 244234 -7386 244854 -7302
rect 244234 -7622 244266 -7386
rect 244502 -7622 244586 -7386
rect 244822 -7622 244854 -7386
rect 244234 -7654 244854 -7622
rect 254194 704838 254814 711590
rect 254194 704602 254226 704838
rect 254462 704602 254546 704838
rect 254782 704602 254814 704838
rect 254194 704518 254814 704602
rect 254194 704282 254226 704518
rect 254462 704282 254546 704518
rect 254782 704282 254814 704518
rect 254194 687854 254814 704282
rect 254194 687618 254226 687854
rect 254462 687618 254546 687854
rect 254782 687618 254814 687854
rect 254194 687534 254814 687618
rect 254194 687298 254226 687534
rect 254462 687298 254546 687534
rect 254782 687298 254814 687534
rect 254194 651854 254814 687298
rect 254194 651618 254226 651854
rect 254462 651618 254546 651854
rect 254782 651618 254814 651854
rect 254194 651534 254814 651618
rect 254194 651298 254226 651534
rect 254462 651298 254546 651534
rect 254782 651298 254814 651534
rect 254194 615854 254814 651298
rect 254194 615618 254226 615854
rect 254462 615618 254546 615854
rect 254782 615618 254814 615854
rect 254194 615534 254814 615618
rect 254194 615298 254226 615534
rect 254462 615298 254546 615534
rect 254782 615298 254814 615534
rect 254194 579854 254814 615298
rect 254194 579618 254226 579854
rect 254462 579618 254546 579854
rect 254782 579618 254814 579854
rect 254194 579534 254814 579618
rect 254194 579298 254226 579534
rect 254462 579298 254546 579534
rect 254782 579298 254814 579534
rect 254194 543854 254814 579298
rect 254194 543618 254226 543854
rect 254462 543618 254546 543854
rect 254782 543618 254814 543854
rect 254194 543534 254814 543618
rect 254194 543298 254226 543534
rect 254462 543298 254546 543534
rect 254782 543298 254814 543534
rect 254194 507854 254814 543298
rect 254194 507618 254226 507854
rect 254462 507618 254546 507854
rect 254782 507618 254814 507854
rect 254194 507534 254814 507618
rect 254194 507298 254226 507534
rect 254462 507298 254546 507534
rect 254782 507298 254814 507534
rect 254194 471854 254814 507298
rect 254194 471618 254226 471854
rect 254462 471618 254546 471854
rect 254782 471618 254814 471854
rect 254194 471534 254814 471618
rect 254194 471298 254226 471534
rect 254462 471298 254546 471534
rect 254782 471298 254814 471534
rect 254194 435854 254814 471298
rect 254194 435618 254226 435854
rect 254462 435618 254546 435854
rect 254782 435618 254814 435854
rect 254194 435534 254814 435618
rect 254194 435298 254226 435534
rect 254462 435298 254546 435534
rect 254782 435298 254814 435534
rect 254194 399854 254814 435298
rect 254194 399618 254226 399854
rect 254462 399618 254546 399854
rect 254782 399618 254814 399854
rect 254194 399534 254814 399618
rect 254194 399298 254226 399534
rect 254462 399298 254546 399534
rect 254782 399298 254814 399534
rect 254194 363854 254814 399298
rect 254194 363618 254226 363854
rect 254462 363618 254546 363854
rect 254782 363618 254814 363854
rect 254194 363534 254814 363618
rect 254194 363298 254226 363534
rect 254462 363298 254546 363534
rect 254782 363298 254814 363534
rect 254194 327854 254814 363298
rect 254194 327618 254226 327854
rect 254462 327618 254546 327854
rect 254782 327618 254814 327854
rect 254194 327534 254814 327618
rect 254194 327298 254226 327534
rect 254462 327298 254546 327534
rect 254782 327298 254814 327534
rect 254194 291854 254814 327298
rect 254194 291618 254226 291854
rect 254462 291618 254546 291854
rect 254782 291618 254814 291854
rect 254194 291534 254814 291618
rect 254194 291298 254226 291534
rect 254462 291298 254546 291534
rect 254782 291298 254814 291534
rect 254194 255854 254814 291298
rect 254194 255618 254226 255854
rect 254462 255618 254546 255854
rect 254782 255618 254814 255854
rect 254194 255534 254814 255618
rect 254194 255298 254226 255534
rect 254462 255298 254546 255534
rect 254782 255298 254814 255534
rect 254194 219854 254814 255298
rect 254194 219618 254226 219854
rect 254462 219618 254546 219854
rect 254782 219618 254814 219854
rect 254194 219534 254814 219618
rect 254194 219298 254226 219534
rect 254462 219298 254546 219534
rect 254782 219298 254814 219534
rect 254194 183854 254814 219298
rect 254194 183618 254226 183854
rect 254462 183618 254546 183854
rect 254782 183618 254814 183854
rect 254194 183534 254814 183618
rect 254194 183298 254226 183534
rect 254462 183298 254546 183534
rect 254782 183298 254814 183534
rect 254194 147854 254814 183298
rect 254194 147618 254226 147854
rect 254462 147618 254546 147854
rect 254782 147618 254814 147854
rect 254194 147534 254814 147618
rect 254194 147298 254226 147534
rect 254462 147298 254546 147534
rect 254782 147298 254814 147534
rect 254194 111854 254814 147298
rect 254194 111618 254226 111854
rect 254462 111618 254546 111854
rect 254782 111618 254814 111854
rect 254194 111534 254814 111618
rect 254194 111298 254226 111534
rect 254462 111298 254546 111534
rect 254782 111298 254814 111534
rect 254194 75854 254814 111298
rect 254194 75618 254226 75854
rect 254462 75618 254546 75854
rect 254782 75618 254814 75854
rect 254194 75534 254814 75618
rect 254194 75298 254226 75534
rect 254462 75298 254546 75534
rect 254782 75298 254814 75534
rect 254194 39854 254814 75298
rect 254194 39618 254226 39854
rect 254462 39618 254546 39854
rect 254782 39618 254814 39854
rect 254194 39534 254814 39618
rect 254194 39298 254226 39534
rect 254462 39298 254546 39534
rect 254782 39298 254814 39534
rect 254194 3854 254814 39298
rect 254194 3618 254226 3854
rect 254462 3618 254546 3854
rect 254782 3618 254814 3854
rect 254194 3534 254814 3618
rect 254194 3298 254226 3534
rect 254462 3298 254546 3534
rect 254782 3298 254814 3534
rect 254194 -346 254814 3298
rect 254194 -582 254226 -346
rect 254462 -582 254546 -346
rect 254782 -582 254814 -346
rect 254194 -666 254814 -582
rect 254194 -902 254226 -666
rect 254462 -902 254546 -666
rect 254782 -902 254814 -666
rect 254194 -7654 254814 -902
rect 257914 705798 258534 711590
rect 257914 705562 257946 705798
rect 258182 705562 258266 705798
rect 258502 705562 258534 705798
rect 257914 705478 258534 705562
rect 257914 705242 257946 705478
rect 258182 705242 258266 705478
rect 258502 705242 258534 705478
rect 257914 691574 258534 705242
rect 257914 691338 257946 691574
rect 258182 691338 258266 691574
rect 258502 691338 258534 691574
rect 257914 691254 258534 691338
rect 257914 691018 257946 691254
rect 258182 691018 258266 691254
rect 258502 691018 258534 691254
rect 257914 655574 258534 691018
rect 257914 655338 257946 655574
rect 258182 655338 258266 655574
rect 258502 655338 258534 655574
rect 257914 655254 258534 655338
rect 257914 655018 257946 655254
rect 258182 655018 258266 655254
rect 258502 655018 258534 655254
rect 257914 619574 258534 655018
rect 257914 619338 257946 619574
rect 258182 619338 258266 619574
rect 258502 619338 258534 619574
rect 257914 619254 258534 619338
rect 257914 619018 257946 619254
rect 258182 619018 258266 619254
rect 258502 619018 258534 619254
rect 257914 583574 258534 619018
rect 257914 583338 257946 583574
rect 258182 583338 258266 583574
rect 258502 583338 258534 583574
rect 257914 583254 258534 583338
rect 257914 583018 257946 583254
rect 258182 583018 258266 583254
rect 258502 583018 258534 583254
rect 257914 547574 258534 583018
rect 257914 547338 257946 547574
rect 258182 547338 258266 547574
rect 258502 547338 258534 547574
rect 257914 547254 258534 547338
rect 257914 547018 257946 547254
rect 258182 547018 258266 547254
rect 258502 547018 258534 547254
rect 257914 511574 258534 547018
rect 257914 511338 257946 511574
rect 258182 511338 258266 511574
rect 258502 511338 258534 511574
rect 257914 511254 258534 511338
rect 257914 511018 257946 511254
rect 258182 511018 258266 511254
rect 258502 511018 258534 511254
rect 257914 475574 258534 511018
rect 257914 475338 257946 475574
rect 258182 475338 258266 475574
rect 258502 475338 258534 475574
rect 257914 475254 258534 475338
rect 257914 475018 257946 475254
rect 258182 475018 258266 475254
rect 258502 475018 258534 475254
rect 257914 439574 258534 475018
rect 257914 439338 257946 439574
rect 258182 439338 258266 439574
rect 258502 439338 258534 439574
rect 257914 439254 258534 439338
rect 257914 439018 257946 439254
rect 258182 439018 258266 439254
rect 258502 439018 258534 439254
rect 257914 403574 258534 439018
rect 257914 403338 257946 403574
rect 258182 403338 258266 403574
rect 258502 403338 258534 403574
rect 257914 403254 258534 403338
rect 257914 403018 257946 403254
rect 258182 403018 258266 403254
rect 258502 403018 258534 403254
rect 257914 367574 258534 403018
rect 257914 367338 257946 367574
rect 258182 367338 258266 367574
rect 258502 367338 258534 367574
rect 257914 367254 258534 367338
rect 257914 367018 257946 367254
rect 258182 367018 258266 367254
rect 258502 367018 258534 367254
rect 257914 331574 258534 367018
rect 257914 331338 257946 331574
rect 258182 331338 258266 331574
rect 258502 331338 258534 331574
rect 257914 331254 258534 331338
rect 257914 331018 257946 331254
rect 258182 331018 258266 331254
rect 258502 331018 258534 331254
rect 257914 295574 258534 331018
rect 257914 295338 257946 295574
rect 258182 295338 258266 295574
rect 258502 295338 258534 295574
rect 257914 295254 258534 295338
rect 257914 295018 257946 295254
rect 258182 295018 258266 295254
rect 258502 295018 258534 295254
rect 257914 259574 258534 295018
rect 257914 259338 257946 259574
rect 258182 259338 258266 259574
rect 258502 259338 258534 259574
rect 257914 259254 258534 259338
rect 257914 259018 257946 259254
rect 258182 259018 258266 259254
rect 258502 259018 258534 259254
rect 257914 223574 258534 259018
rect 257914 223338 257946 223574
rect 258182 223338 258266 223574
rect 258502 223338 258534 223574
rect 257914 223254 258534 223338
rect 257914 223018 257946 223254
rect 258182 223018 258266 223254
rect 258502 223018 258534 223254
rect 257914 187574 258534 223018
rect 257914 187338 257946 187574
rect 258182 187338 258266 187574
rect 258502 187338 258534 187574
rect 257914 187254 258534 187338
rect 257914 187018 257946 187254
rect 258182 187018 258266 187254
rect 258502 187018 258534 187254
rect 257914 151574 258534 187018
rect 257914 151338 257946 151574
rect 258182 151338 258266 151574
rect 258502 151338 258534 151574
rect 257914 151254 258534 151338
rect 257914 151018 257946 151254
rect 258182 151018 258266 151254
rect 258502 151018 258534 151254
rect 257914 115574 258534 151018
rect 257914 115338 257946 115574
rect 258182 115338 258266 115574
rect 258502 115338 258534 115574
rect 257914 115254 258534 115338
rect 257914 115018 257946 115254
rect 258182 115018 258266 115254
rect 258502 115018 258534 115254
rect 257914 79574 258534 115018
rect 257914 79338 257946 79574
rect 258182 79338 258266 79574
rect 258502 79338 258534 79574
rect 257914 79254 258534 79338
rect 257914 79018 257946 79254
rect 258182 79018 258266 79254
rect 258502 79018 258534 79254
rect 257914 43574 258534 79018
rect 257914 43338 257946 43574
rect 258182 43338 258266 43574
rect 258502 43338 258534 43574
rect 257914 43254 258534 43338
rect 257914 43018 257946 43254
rect 258182 43018 258266 43254
rect 258502 43018 258534 43254
rect 257914 7574 258534 43018
rect 257914 7338 257946 7574
rect 258182 7338 258266 7574
rect 258502 7338 258534 7574
rect 257914 7254 258534 7338
rect 257914 7018 257946 7254
rect 258182 7018 258266 7254
rect 258502 7018 258534 7254
rect 257914 -1306 258534 7018
rect 257914 -1542 257946 -1306
rect 258182 -1542 258266 -1306
rect 258502 -1542 258534 -1306
rect 257914 -1626 258534 -1542
rect 257914 -1862 257946 -1626
rect 258182 -1862 258266 -1626
rect 258502 -1862 258534 -1626
rect 257914 -7654 258534 -1862
rect 261634 706758 262254 711590
rect 261634 706522 261666 706758
rect 261902 706522 261986 706758
rect 262222 706522 262254 706758
rect 261634 706438 262254 706522
rect 261634 706202 261666 706438
rect 261902 706202 261986 706438
rect 262222 706202 262254 706438
rect 261634 695294 262254 706202
rect 261634 695058 261666 695294
rect 261902 695058 261986 695294
rect 262222 695058 262254 695294
rect 261634 694974 262254 695058
rect 261634 694738 261666 694974
rect 261902 694738 261986 694974
rect 262222 694738 262254 694974
rect 261634 659294 262254 694738
rect 261634 659058 261666 659294
rect 261902 659058 261986 659294
rect 262222 659058 262254 659294
rect 261634 658974 262254 659058
rect 261634 658738 261666 658974
rect 261902 658738 261986 658974
rect 262222 658738 262254 658974
rect 261634 623294 262254 658738
rect 261634 623058 261666 623294
rect 261902 623058 261986 623294
rect 262222 623058 262254 623294
rect 261634 622974 262254 623058
rect 261634 622738 261666 622974
rect 261902 622738 261986 622974
rect 262222 622738 262254 622974
rect 261634 587294 262254 622738
rect 261634 587058 261666 587294
rect 261902 587058 261986 587294
rect 262222 587058 262254 587294
rect 261634 586974 262254 587058
rect 261634 586738 261666 586974
rect 261902 586738 261986 586974
rect 262222 586738 262254 586974
rect 261634 551294 262254 586738
rect 261634 551058 261666 551294
rect 261902 551058 261986 551294
rect 262222 551058 262254 551294
rect 261634 550974 262254 551058
rect 261634 550738 261666 550974
rect 261902 550738 261986 550974
rect 262222 550738 262254 550974
rect 261634 515294 262254 550738
rect 261634 515058 261666 515294
rect 261902 515058 261986 515294
rect 262222 515058 262254 515294
rect 261634 514974 262254 515058
rect 261634 514738 261666 514974
rect 261902 514738 261986 514974
rect 262222 514738 262254 514974
rect 261634 479294 262254 514738
rect 261634 479058 261666 479294
rect 261902 479058 261986 479294
rect 262222 479058 262254 479294
rect 261634 478974 262254 479058
rect 261634 478738 261666 478974
rect 261902 478738 261986 478974
rect 262222 478738 262254 478974
rect 261634 443294 262254 478738
rect 261634 443058 261666 443294
rect 261902 443058 261986 443294
rect 262222 443058 262254 443294
rect 261634 442974 262254 443058
rect 261634 442738 261666 442974
rect 261902 442738 261986 442974
rect 262222 442738 262254 442974
rect 261634 407294 262254 442738
rect 261634 407058 261666 407294
rect 261902 407058 261986 407294
rect 262222 407058 262254 407294
rect 261634 406974 262254 407058
rect 261634 406738 261666 406974
rect 261902 406738 261986 406974
rect 262222 406738 262254 406974
rect 261634 371294 262254 406738
rect 261634 371058 261666 371294
rect 261902 371058 261986 371294
rect 262222 371058 262254 371294
rect 261634 370974 262254 371058
rect 261634 370738 261666 370974
rect 261902 370738 261986 370974
rect 262222 370738 262254 370974
rect 261634 335294 262254 370738
rect 261634 335058 261666 335294
rect 261902 335058 261986 335294
rect 262222 335058 262254 335294
rect 261634 334974 262254 335058
rect 261634 334738 261666 334974
rect 261902 334738 261986 334974
rect 262222 334738 262254 334974
rect 261634 299294 262254 334738
rect 261634 299058 261666 299294
rect 261902 299058 261986 299294
rect 262222 299058 262254 299294
rect 261634 298974 262254 299058
rect 261634 298738 261666 298974
rect 261902 298738 261986 298974
rect 262222 298738 262254 298974
rect 261634 263294 262254 298738
rect 261634 263058 261666 263294
rect 261902 263058 261986 263294
rect 262222 263058 262254 263294
rect 261634 262974 262254 263058
rect 261634 262738 261666 262974
rect 261902 262738 261986 262974
rect 262222 262738 262254 262974
rect 261634 227294 262254 262738
rect 261634 227058 261666 227294
rect 261902 227058 261986 227294
rect 262222 227058 262254 227294
rect 261634 226974 262254 227058
rect 261634 226738 261666 226974
rect 261902 226738 261986 226974
rect 262222 226738 262254 226974
rect 261634 191294 262254 226738
rect 261634 191058 261666 191294
rect 261902 191058 261986 191294
rect 262222 191058 262254 191294
rect 261634 190974 262254 191058
rect 261634 190738 261666 190974
rect 261902 190738 261986 190974
rect 262222 190738 262254 190974
rect 261634 155294 262254 190738
rect 261634 155058 261666 155294
rect 261902 155058 261986 155294
rect 262222 155058 262254 155294
rect 261634 154974 262254 155058
rect 261634 154738 261666 154974
rect 261902 154738 261986 154974
rect 262222 154738 262254 154974
rect 261634 119294 262254 154738
rect 261634 119058 261666 119294
rect 261902 119058 261986 119294
rect 262222 119058 262254 119294
rect 261634 118974 262254 119058
rect 261634 118738 261666 118974
rect 261902 118738 261986 118974
rect 262222 118738 262254 118974
rect 261634 83294 262254 118738
rect 261634 83058 261666 83294
rect 261902 83058 261986 83294
rect 262222 83058 262254 83294
rect 261634 82974 262254 83058
rect 261634 82738 261666 82974
rect 261902 82738 261986 82974
rect 262222 82738 262254 82974
rect 261634 47294 262254 82738
rect 261634 47058 261666 47294
rect 261902 47058 261986 47294
rect 262222 47058 262254 47294
rect 261634 46974 262254 47058
rect 261634 46738 261666 46974
rect 261902 46738 261986 46974
rect 262222 46738 262254 46974
rect 261634 11294 262254 46738
rect 261634 11058 261666 11294
rect 261902 11058 261986 11294
rect 262222 11058 262254 11294
rect 261634 10974 262254 11058
rect 261634 10738 261666 10974
rect 261902 10738 261986 10974
rect 262222 10738 262254 10974
rect 261634 -2266 262254 10738
rect 261634 -2502 261666 -2266
rect 261902 -2502 261986 -2266
rect 262222 -2502 262254 -2266
rect 261634 -2586 262254 -2502
rect 261634 -2822 261666 -2586
rect 261902 -2822 261986 -2586
rect 262222 -2822 262254 -2586
rect 261634 -7654 262254 -2822
rect 265354 707718 265974 711590
rect 265354 707482 265386 707718
rect 265622 707482 265706 707718
rect 265942 707482 265974 707718
rect 265354 707398 265974 707482
rect 265354 707162 265386 707398
rect 265622 707162 265706 707398
rect 265942 707162 265974 707398
rect 265354 699014 265974 707162
rect 265354 698778 265386 699014
rect 265622 698778 265706 699014
rect 265942 698778 265974 699014
rect 265354 698694 265974 698778
rect 265354 698458 265386 698694
rect 265622 698458 265706 698694
rect 265942 698458 265974 698694
rect 265354 663014 265974 698458
rect 265354 662778 265386 663014
rect 265622 662778 265706 663014
rect 265942 662778 265974 663014
rect 265354 662694 265974 662778
rect 265354 662458 265386 662694
rect 265622 662458 265706 662694
rect 265942 662458 265974 662694
rect 265354 627014 265974 662458
rect 265354 626778 265386 627014
rect 265622 626778 265706 627014
rect 265942 626778 265974 627014
rect 265354 626694 265974 626778
rect 265354 626458 265386 626694
rect 265622 626458 265706 626694
rect 265942 626458 265974 626694
rect 265354 591014 265974 626458
rect 265354 590778 265386 591014
rect 265622 590778 265706 591014
rect 265942 590778 265974 591014
rect 265354 590694 265974 590778
rect 265354 590458 265386 590694
rect 265622 590458 265706 590694
rect 265942 590458 265974 590694
rect 265354 555014 265974 590458
rect 265354 554778 265386 555014
rect 265622 554778 265706 555014
rect 265942 554778 265974 555014
rect 265354 554694 265974 554778
rect 265354 554458 265386 554694
rect 265622 554458 265706 554694
rect 265942 554458 265974 554694
rect 265354 519014 265974 554458
rect 265354 518778 265386 519014
rect 265622 518778 265706 519014
rect 265942 518778 265974 519014
rect 265354 518694 265974 518778
rect 265354 518458 265386 518694
rect 265622 518458 265706 518694
rect 265942 518458 265974 518694
rect 265354 483014 265974 518458
rect 265354 482778 265386 483014
rect 265622 482778 265706 483014
rect 265942 482778 265974 483014
rect 265354 482694 265974 482778
rect 265354 482458 265386 482694
rect 265622 482458 265706 482694
rect 265942 482458 265974 482694
rect 265354 447014 265974 482458
rect 265354 446778 265386 447014
rect 265622 446778 265706 447014
rect 265942 446778 265974 447014
rect 265354 446694 265974 446778
rect 265354 446458 265386 446694
rect 265622 446458 265706 446694
rect 265942 446458 265974 446694
rect 265354 411014 265974 446458
rect 265354 410778 265386 411014
rect 265622 410778 265706 411014
rect 265942 410778 265974 411014
rect 265354 410694 265974 410778
rect 265354 410458 265386 410694
rect 265622 410458 265706 410694
rect 265942 410458 265974 410694
rect 265354 375014 265974 410458
rect 265354 374778 265386 375014
rect 265622 374778 265706 375014
rect 265942 374778 265974 375014
rect 265354 374694 265974 374778
rect 265354 374458 265386 374694
rect 265622 374458 265706 374694
rect 265942 374458 265974 374694
rect 265354 339014 265974 374458
rect 265354 338778 265386 339014
rect 265622 338778 265706 339014
rect 265942 338778 265974 339014
rect 265354 338694 265974 338778
rect 265354 338458 265386 338694
rect 265622 338458 265706 338694
rect 265942 338458 265974 338694
rect 265354 303014 265974 338458
rect 265354 302778 265386 303014
rect 265622 302778 265706 303014
rect 265942 302778 265974 303014
rect 265354 302694 265974 302778
rect 265354 302458 265386 302694
rect 265622 302458 265706 302694
rect 265942 302458 265974 302694
rect 265354 267014 265974 302458
rect 265354 266778 265386 267014
rect 265622 266778 265706 267014
rect 265942 266778 265974 267014
rect 265354 266694 265974 266778
rect 265354 266458 265386 266694
rect 265622 266458 265706 266694
rect 265942 266458 265974 266694
rect 265354 231014 265974 266458
rect 265354 230778 265386 231014
rect 265622 230778 265706 231014
rect 265942 230778 265974 231014
rect 265354 230694 265974 230778
rect 265354 230458 265386 230694
rect 265622 230458 265706 230694
rect 265942 230458 265974 230694
rect 265354 195014 265974 230458
rect 265354 194778 265386 195014
rect 265622 194778 265706 195014
rect 265942 194778 265974 195014
rect 265354 194694 265974 194778
rect 265354 194458 265386 194694
rect 265622 194458 265706 194694
rect 265942 194458 265974 194694
rect 265354 159014 265974 194458
rect 265354 158778 265386 159014
rect 265622 158778 265706 159014
rect 265942 158778 265974 159014
rect 265354 158694 265974 158778
rect 265354 158458 265386 158694
rect 265622 158458 265706 158694
rect 265942 158458 265974 158694
rect 265354 123014 265974 158458
rect 265354 122778 265386 123014
rect 265622 122778 265706 123014
rect 265942 122778 265974 123014
rect 265354 122694 265974 122778
rect 265354 122458 265386 122694
rect 265622 122458 265706 122694
rect 265942 122458 265974 122694
rect 265354 87014 265974 122458
rect 265354 86778 265386 87014
rect 265622 86778 265706 87014
rect 265942 86778 265974 87014
rect 265354 86694 265974 86778
rect 265354 86458 265386 86694
rect 265622 86458 265706 86694
rect 265942 86458 265974 86694
rect 265354 51014 265974 86458
rect 265354 50778 265386 51014
rect 265622 50778 265706 51014
rect 265942 50778 265974 51014
rect 265354 50694 265974 50778
rect 265354 50458 265386 50694
rect 265622 50458 265706 50694
rect 265942 50458 265974 50694
rect 265354 15014 265974 50458
rect 265354 14778 265386 15014
rect 265622 14778 265706 15014
rect 265942 14778 265974 15014
rect 265354 14694 265974 14778
rect 265354 14458 265386 14694
rect 265622 14458 265706 14694
rect 265942 14458 265974 14694
rect 265354 -3226 265974 14458
rect 265354 -3462 265386 -3226
rect 265622 -3462 265706 -3226
rect 265942 -3462 265974 -3226
rect 265354 -3546 265974 -3462
rect 265354 -3782 265386 -3546
rect 265622 -3782 265706 -3546
rect 265942 -3782 265974 -3546
rect 265354 -7654 265974 -3782
rect 269074 708678 269694 711590
rect 269074 708442 269106 708678
rect 269342 708442 269426 708678
rect 269662 708442 269694 708678
rect 269074 708358 269694 708442
rect 269074 708122 269106 708358
rect 269342 708122 269426 708358
rect 269662 708122 269694 708358
rect 269074 666734 269694 708122
rect 269074 666498 269106 666734
rect 269342 666498 269426 666734
rect 269662 666498 269694 666734
rect 269074 666414 269694 666498
rect 269074 666178 269106 666414
rect 269342 666178 269426 666414
rect 269662 666178 269694 666414
rect 269074 630734 269694 666178
rect 269074 630498 269106 630734
rect 269342 630498 269426 630734
rect 269662 630498 269694 630734
rect 269074 630414 269694 630498
rect 269074 630178 269106 630414
rect 269342 630178 269426 630414
rect 269662 630178 269694 630414
rect 269074 594734 269694 630178
rect 269074 594498 269106 594734
rect 269342 594498 269426 594734
rect 269662 594498 269694 594734
rect 269074 594414 269694 594498
rect 269074 594178 269106 594414
rect 269342 594178 269426 594414
rect 269662 594178 269694 594414
rect 269074 558734 269694 594178
rect 269074 558498 269106 558734
rect 269342 558498 269426 558734
rect 269662 558498 269694 558734
rect 269074 558414 269694 558498
rect 269074 558178 269106 558414
rect 269342 558178 269426 558414
rect 269662 558178 269694 558414
rect 269074 522734 269694 558178
rect 269074 522498 269106 522734
rect 269342 522498 269426 522734
rect 269662 522498 269694 522734
rect 269074 522414 269694 522498
rect 269074 522178 269106 522414
rect 269342 522178 269426 522414
rect 269662 522178 269694 522414
rect 269074 486734 269694 522178
rect 269074 486498 269106 486734
rect 269342 486498 269426 486734
rect 269662 486498 269694 486734
rect 269074 486414 269694 486498
rect 269074 486178 269106 486414
rect 269342 486178 269426 486414
rect 269662 486178 269694 486414
rect 269074 450734 269694 486178
rect 269074 450498 269106 450734
rect 269342 450498 269426 450734
rect 269662 450498 269694 450734
rect 269074 450414 269694 450498
rect 269074 450178 269106 450414
rect 269342 450178 269426 450414
rect 269662 450178 269694 450414
rect 269074 414734 269694 450178
rect 269074 414498 269106 414734
rect 269342 414498 269426 414734
rect 269662 414498 269694 414734
rect 269074 414414 269694 414498
rect 269074 414178 269106 414414
rect 269342 414178 269426 414414
rect 269662 414178 269694 414414
rect 269074 378734 269694 414178
rect 269074 378498 269106 378734
rect 269342 378498 269426 378734
rect 269662 378498 269694 378734
rect 269074 378414 269694 378498
rect 269074 378178 269106 378414
rect 269342 378178 269426 378414
rect 269662 378178 269694 378414
rect 269074 342734 269694 378178
rect 269074 342498 269106 342734
rect 269342 342498 269426 342734
rect 269662 342498 269694 342734
rect 269074 342414 269694 342498
rect 269074 342178 269106 342414
rect 269342 342178 269426 342414
rect 269662 342178 269694 342414
rect 269074 306734 269694 342178
rect 269074 306498 269106 306734
rect 269342 306498 269426 306734
rect 269662 306498 269694 306734
rect 269074 306414 269694 306498
rect 269074 306178 269106 306414
rect 269342 306178 269426 306414
rect 269662 306178 269694 306414
rect 269074 270734 269694 306178
rect 269074 270498 269106 270734
rect 269342 270498 269426 270734
rect 269662 270498 269694 270734
rect 269074 270414 269694 270498
rect 269074 270178 269106 270414
rect 269342 270178 269426 270414
rect 269662 270178 269694 270414
rect 269074 234734 269694 270178
rect 269074 234498 269106 234734
rect 269342 234498 269426 234734
rect 269662 234498 269694 234734
rect 269074 234414 269694 234498
rect 269074 234178 269106 234414
rect 269342 234178 269426 234414
rect 269662 234178 269694 234414
rect 269074 198734 269694 234178
rect 269074 198498 269106 198734
rect 269342 198498 269426 198734
rect 269662 198498 269694 198734
rect 269074 198414 269694 198498
rect 269074 198178 269106 198414
rect 269342 198178 269426 198414
rect 269662 198178 269694 198414
rect 269074 162734 269694 198178
rect 269074 162498 269106 162734
rect 269342 162498 269426 162734
rect 269662 162498 269694 162734
rect 269074 162414 269694 162498
rect 269074 162178 269106 162414
rect 269342 162178 269426 162414
rect 269662 162178 269694 162414
rect 269074 126734 269694 162178
rect 269074 126498 269106 126734
rect 269342 126498 269426 126734
rect 269662 126498 269694 126734
rect 269074 126414 269694 126498
rect 269074 126178 269106 126414
rect 269342 126178 269426 126414
rect 269662 126178 269694 126414
rect 269074 90734 269694 126178
rect 269074 90498 269106 90734
rect 269342 90498 269426 90734
rect 269662 90498 269694 90734
rect 269074 90414 269694 90498
rect 269074 90178 269106 90414
rect 269342 90178 269426 90414
rect 269662 90178 269694 90414
rect 269074 54734 269694 90178
rect 269074 54498 269106 54734
rect 269342 54498 269426 54734
rect 269662 54498 269694 54734
rect 269074 54414 269694 54498
rect 269074 54178 269106 54414
rect 269342 54178 269426 54414
rect 269662 54178 269694 54414
rect 269074 18734 269694 54178
rect 269074 18498 269106 18734
rect 269342 18498 269426 18734
rect 269662 18498 269694 18734
rect 269074 18414 269694 18498
rect 269074 18178 269106 18414
rect 269342 18178 269426 18414
rect 269662 18178 269694 18414
rect 269074 -4186 269694 18178
rect 269074 -4422 269106 -4186
rect 269342 -4422 269426 -4186
rect 269662 -4422 269694 -4186
rect 269074 -4506 269694 -4422
rect 269074 -4742 269106 -4506
rect 269342 -4742 269426 -4506
rect 269662 -4742 269694 -4506
rect 269074 -7654 269694 -4742
rect 272794 709638 273414 711590
rect 272794 709402 272826 709638
rect 273062 709402 273146 709638
rect 273382 709402 273414 709638
rect 272794 709318 273414 709402
rect 272794 709082 272826 709318
rect 273062 709082 273146 709318
rect 273382 709082 273414 709318
rect 272794 670454 273414 709082
rect 272794 670218 272826 670454
rect 273062 670218 273146 670454
rect 273382 670218 273414 670454
rect 272794 670134 273414 670218
rect 272794 669898 272826 670134
rect 273062 669898 273146 670134
rect 273382 669898 273414 670134
rect 272794 634454 273414 669898
rect 272794 634218 272826 634454
rect 273062 634218 273146 634454
rect 273382 634218 273414 634454
rect 272794 634134 273414 634218
rect 272794 633898 272826 634134
rect 273062 633898 273146 634134
rect 273382 633898 273414 634134
rect 272794 598454 273414 633898
rect 272794 598218 272826 598454
rect 273062 598218 273146 598454
rect 273382 598218 273414 598454
rect 272794 598134 273414 598218
rect 272794 597898 272826 598134
rect 273062 597898 273146 598134
rect 273382 597898 273414 598134
rect 272794 562454 273414 597898
rect 272794 562218 272826 562454
rect 273062 562218 273146 562454
rect 273382 562218 273414 562454
rect 272794 562134 273414 562218
rect 272794 561898 272826 562134
rect 273062 561898 273146 562134
rect 273382 561898 273414 562134
rect 272794 526454 273414 561898
rect 272794 526218 272826 526454
rect 273062 526218 273146 526454
rect 273382 526218 273414 526454
rect 272794 526134 273414 526218
rect 272794 525898 272826 526134
rect 273062 525898 273146 526134
rect 273382 525898 273414 526134
rect 272794 490454 273414 525898
rect 272794 490218 272826 490454
rect 273062 490218 273146 490454
rect 273382 490218 273414 490454
rect 272794 490134 273414 490218
rect 272794 489898 272826 490134
rect 273062 489898 273146 490134
rect 273382 489898 273414 490134
rect 272794 454454 273414 489898
rect 272794 454218 272826 454454
rect 273062 454218 273146 454454
rect 273382 454218 273414 454454
rect 272794 454134 273414 454218
rect 272794 453898 272826 454134
rect 273062 453898 273146 454134
rect 273382 453898 273414 454134
rect 272794 418454 273414 453898
rect 272794 418218 272826 418454
rect 273062 418218 273146 418454
rect 273382 418218 273414 418454
rect 272794 418134 273414 418218
rect 272794 417898 272826 418134
rect 273062 417898 273146 418134
rect 273382 417898 273414 418134
rect 272794 382454 273414 417898
rect 272794 382218 272826 382454
rect 273062 382218 273146 382454
rect 273382 382218 273414 382454
rect 272794 382134 273414 382218
rect 272794 381898 272826 382134
rect 273062 381898 273146 382134
rect 273382 381898 273414 382134
rect 272794 346454 273414 381898
rect 272794 346218 272826 346454
rect 273062 346218 273146 346454
rect 273382 346218 273414 346454
rect 272794 346134 273414 346218
rect 272794 345898 272826 346134
rect 273062 345898 273146 346134
rect 273382 345898 273414 346134
rect 272794 310454 273414 345898
rect 272794 310218 272826 310454
rect 273062 310218 273146 310454
rect 273382 310218 273414 310454
rect 272794 310134 273414 310218
rect 272794 309898 272826 310134
rect 273062 309898 273146 310134
rect 273382 309898 273414 310134
rect 272794 274454 273414 309898
rect 272794 274218 272826 274454
rect 273062 274218 273146 274454
rect 273382 274218 273414 274454
rect 272794 274134 273414 274218
rect 272794 273898 272826 274134
rect 273062 273898 273146 274134
rect 273382 273898 273414 274134
rect 272794 238454 273414 273898
rect 272794 238218 272826 238454
rect 273062 238218 273146 238454
rect 273382 238218 273414 238454
rect 272794 238134 273414 238218
rect 272794 237898 272826 238134
rect 273062 237898 273146 238134
rect 273382 237898 273414 238134
rect 272794 202454 273414 237898
rect 272794 202218 272826 202454
rect 273062 202218 273146 202454
rect 273382 202218 273414 202454
rect 272794 202134 273414 202218
rect 272794 201898 272826 202134
rect 273062 201898 273146 202134
rect 273382 201898 273414 202134
rect 272794 166454 273414 201898
rect 272794 166218 272826 166454
rect 273062 166218 273146 166454
rect 273382 166218 273414 166454
rect 272794 166134 273414 166218
rect 272794 165898 272826 166134
rect 273062 165898 273146 166134
rect 273382 165898 273414 166134
rect 272794 130454 273414 165898
rect 272794 130218 272826 130454
rect 273062 130218 273146 130454
rect 273382 130218 273414 130454
rect 272794 130134 273414 130218
rect 272794 129898 272826 130134
rect 273062 129898 273146 130134
rect 273382 129898 273414 130134
rect 272794 94454 273414 129898
rect 272794 94218 272826 94454
rect 273062 94218 273146 94454
rect 273382 94218 273414 94454
rect 272794 94134 273414 94218
rect 272794 93898 272826 94134
rect 273062 93898 273146 94134
rect 273382 93898 273414 94134
rect 272794 58454 273414 93898
rect 272794 58218 272826 58454
rect 273062 58218 273146 58454
rect 273382 58218 273414 58454
rect 272794 58134 273414 58218
rect 272794 57898 272826 58134
rect 273062 57898 273146 58134
rect 273382 57898 273414 58134
rect 272794 22454 273414 57898
rect 272794 22218 272826 22454
rect 273062 22218 273146 22454
rect 273382 22218 273414 22454
rect 272794 22134 273414 22218
rect 272794 21898 272826 22134
rect 273062 21898 273146 22134
rect 273382 21898 273414 22134
rect 272794 -5146 273414 21898
rect 272794 -5382 272826 -5146
rect 273062 -5382 273146 -5146
rect 273382 -5382 273414 -5146
rect 272794 -5466 273414 -5382
rect 272794 -5702 272826 -5466
rect 273062 -5702 273146 -5466
rect 273382 -5702 273414 -5466
rect 272794 -7654 273414 -5702
rect 276514 710598 277134 711590
rect 276514 710362 276546 710598
rect 276782 710362 276866 710598
rect 277102 710362 277134 710598
rect 276514 710278 277134 710362
rect 276514 710042 276546 710278
rect 276782 710042 276866 710278
rect 277102 710042 277134 710278
rect 276514 674174 277134 710042
rect 276514 673938 276546 674174
rect 276782 673938 276866 674174
rect 277102 673938 277134 674174
rect 276514 673854 277134 673938
rect 276514 673618 276546 673854
rect 276782 673618 276866 673854
rect 277102 673618 277134 673854
rect 276514 638174 277134 673618
rect 276514 637938 276546 638174
rect 276782 637938 276866 638174
rect 277102 637938 277134 638174
rect 276514 637854 277134 637938
rect 276514 637618 276546 637854
rect 276782 637618 276866 637854
rect 277102 637618 277134 637854
rect 276514 602174 277134 637618
rect 276514 601938 276546 602174
rect 276782 601938 276866 602174
rect 277102 601938 277134 602174
rect 276514 601854 277134 601938
rect 276514 601618 276546 601854
rect 276782 601618 276866 601854
rect 277102 601618 277134 601854
rect 276514 566174 277134 601618
rect 276514 565938 276546 566174
rect 276782 565938 276866 566174
rect 277102 565938 277134 566174
rect 276514 565854 277134 565938
rect 276514 565618 276546 565854
rect 276782 565618 276866 565854
rect 277102 565618 277134 565854
rect 276514 530174 277134 565618
rect 276514 529938 276546 530174
rect 276782 529938 276866 530174
rect 277102 529938 277134 530174
rect 276514 529854 277134 529938
rect 276514 529618 276546 529854
rect 276782 529618 276866 529854
rect 277102 529618 277134 529854
rect 276514 494174 277134 529618
rect 276514 493938 276546 494174
rect 276782 493938 276866 494174
rect 277102 493938 277134 494174
rect 276514 493854 277134 493938
rect 276514 493618 276546 493854
rect 276782 493618 276866 493854
rect 277102 493618 277134 493854
rect 276514 458174 277134 493618
rect 276514 457938 276546 458174
rect 276782 457938 276866 458174
rect 277102 457938 277134 458174
rect 276514 457854 277134 457938
rect 276514 457618 276546 457854
rect 276782 457618 276866 457854
rect 277102 457618 277134 457854
rect 276514 422174 277134 457618
rect 276514 421938 276546 422174
rect 276782 421938 276866 422174
rect 277102 421938 277134 422174
rect 276514 421854 277134 421938
rect 276514 421618 276546 421854
rect 276782 421618 276866 421854
rect 277102 421618 277134 421854
rect 276514 386174 277134 421618
rect 276514 385938 276546 386174
rect 276782 385938 276866 386174
rect 277102 385938 277134 386174
rect 276514 385854 277134 385938
rect 276514 385618 276546 385854
rect 276782 385618 276866 385854
rect 277102 385618 277134 385854
rect 276514 350174 277134 385618
rect 276514 349938 276546 350174
rect 276782 349938 276866 350174
rect 277102 349938 277134 350174
rect 276514 349854 277134 349938
rect 276514 349618 276546 349854
rect 276782 349618 276866 349854
rect 277102 349618 277134 349854
rect 276514 314174 277134 349618
rect 276514 313938 276546 314174
rect 276782 313938 276866 314174
rect 277102 313938 277134 314174
rect 276514 313854 277134 313938
rect 276514 313618 276546 313854
rect 276782 313618 276866 313854
rect 277102 313618 277134 313854
rect 276514 278174 277134 313618
rect 276514 277938 276546 278174
rect 276782 277938 276866 278174
rect 277102 277938 277134 278174
rect 276514 277854 277134 277938
rect 276514 277618 276546 277854
rect 276782 277618 276866 277854
rect 277102 277618 277134 277854
rect 276514 242174 277134 277618
rect 276514 241938 276546 242174
rect 276782 241938 276866 242174
rect 277102 241938 277134 242174
rect 276514 241854 277134 241938
rect 276514 241618 276546 241854
rect 276782 241618 276866 241854
rect 277102 241618 277134 241854
rect 276514 206174 277134 241618
rect 276514 205938 276546 206174
rect 276782 205938 276866 206174
rect 277102 205938 277134 206174
rect 276514 205854 277134 205938
rect 276514 205618 276546 205854
rect 276782 205618 276866 205854
rect 277102 205618 277134 205854
rect 276514 170174 277134 205618
rect 276514 169938 276546 170174
rect 276782 169938 276866 170174
rect 277102 169938 277134 170174
rect 276514 169854 277134 169938
rect 276514 169618 276546 169854
rect 276782 169618 276866 169854
rect 277102 169618 277134 169854
rect 276514 134174 277134 169618
rect 276514 133938 276546 134174
rect 276782 133938 276866 134174
rect 277102 133938 277134 134174
rect 276514 133854 277134 133938
rect 276514 133618 276546 133854
rect 276782 133618 276866 133854
rect 277102 133618 277134 133854
rect 276514 98174 277134 133618
rect 276514 97938 276546 98174
rect 276782 97938 276866 98174
rect 277102 97938 277134 98174
rect 276514 97854 277134 97938
rect 276514 97618 276546 97854
rect 276782 97618 276866 97854
rect 277102 97618 277134 97854
rect 276514 62174 277134 97618
rect 276514 61938 276546 62174
rect 276782 61938 276866 62174
rect 277102 61938 277134 62174
rect 276514 61854 277134 61938
rect 276514 61618 276546 61854
rect 276782 61618 276866 61854
rect 277102 61618 277134 61854
rect 276514 26174 277134 61618
rect 276514 25938 276546 26174
rect 276782 25938 276866 26174
rect 277102 25938 277134 26174
rect 276514 25854 277134 25938
rect 276514 25618 276546 25854
rect 276782 25618 276866 25854
rect 277102 25618 277134 25854
rect 276514 -6106 277134 25618
rect 276514 -6342 276546 -6106
rect 276782 -6342 276866 -6106
rect 277102 -6342 277134 -6106
rect 276514 -6426 277134 -6342
rect 276514 -6662 276546 -6426
rect 276782 -6662 276866 -6426
rect 277102 -6662 277134 -6426
rect 276514 -7654 277134 -6662
rect 280234 711558 280854 711590
rect 280234 711322 280266 711558
rect 280502 711322 280586 711558
rect 280822 711322 280854 711558
rect 280234 711238 280854 711322
rect 280234 711002 280266 711238
rect 280502 711002 280586 711238
rect 280822 711002 280854 711238
rect 280234 677894 280854 711002
rect 280234 677658 280266 677894
rect 280502 677658 280586 677894
rect 280822 677658 280854 677894
rect 280234 677574 280854 677658
rect 280234 677338 280266 677574
rect 280502 677338 280586 677574
rect 280822 677338 280854 677574
rect 280234 641894 280854 677338
rect 280234 641658 280266 641894
rect 280502 641658 280586 641894
rect 280822 641658 280854 641894
rect 280234 641574 280854 641658
rect 280234 641338 280266 641574
rect 280502 641338 280586 641574
rect 280822 641338 280854 641574
rect 280234 605894 280854 641338
rect 280234 605658 280266 605894
rect 280502 605658 280586 605894
rect 280822 605658 280854 605894
rect 280234 605574 280854 605658
rect 280234 605338 280266 605574
rect 280502 605338 280586 605574
rect 280822 605338 280854 605574
rect 280234 569894 280854 605338
rect 280234 569658 280266 569894
rect 280502 569658 280586 569894
rect 280822 569658 280854 569894
rect 280234 569574 280854 569658
rect 280234 569338 280266 569574
rect 280502 569338 280586 569574
rect 280822 569338 280854 569574
rect 280234 533894 280854 569338
rect 280234 533658 280266 533894
rect 280502 533658 280586 533894
rect 280822 533658 280854 533894
rect 280234 533574 280854 533658
rect 280234 533338 280266 533574
rect 280502 533338 280586 533574
rect 280822 533338 280854 533574
rect 280234 497894 280854 533338
rect 280234 497658 280266 497894
rect 280502 497658 280586 497894
rect 280822 497658 280854 497894
rect 280234 497574 280854 497658
rect 280234 497338 280266 497574
rect 280502 497338 280586 497574
rect 280822 497338 280854 497574
rect 280234 461894 280854 497338
rect 280234 461658 280266 461894
rect 280502 461658 280586 461894
rect 280822 461658 280854 461894
rect 280234 461574 280854 461658
rect 280234 461338 280266 461574
rect 280502 461338 280586 461574
rect 280822 461338 280854 461574
rect 280234 425894 280854 461338
rect 280234 425658 280266 425894
rect 280502 425658 280586 425894
rect 280822 425658 280854 425894
rect 280234 425574 280854 425658
rect 280234 425338 280266 425574
rect 280502 425338 280586 425574
rect 280822 425338 280854 425574
rect 280234 389894 280854 425338
rect 280234 389658 280266 389894
rect 280502 389658 280586 389894
rect 280822 389658 280854 389894
rect 280234 389574 280854 389658
rect 280234 389338 280266 389574
rect 280502 389338 280586 389574
rect 280822 389338 280854 389574
rect 280234 353894 280854 389338
rect 280234 353658 280266 353894
rect 280502 353658 280586 353894
rect 280822 353658 280854 353894
rect 280234 353574 280854 353658
rect 280234 353338 280266 353574
rect 280502 353338 280586 353574
rect 280822 353338 280854 353574
rect 280234 317894 280854 353338
rect 280234 317658 280266 317894
rect 280502 317658 280586 317894
rect 280822 317658 280854 317894
rect 280234 317574 280854 317658
rect 280234 317338 280266 317574
rect 280502 317338 280586 317574
rect 280822 317338 280854 317574
rect 280234 281894 280854 317338
rect 280234 281658 280266 281894
rect 280502 281658 280586 281894
rect 280822 281658 280854 281894
rect 280234 281574 280854 281658
rect 280234 281338 280266 281574
rect 280502 281338 280586 281574
rect 280822 281338 280854 281574
rect 280234 245894 280854 281338
rect 280234 245658 280266 245894
rect 280502 245658 280586 245894
rect 280822 245658 280854 245894
rect 280234 245574 280854 245658
rect 280234 245338 280266 245574
rect 280502 245338 280586 245574
rect 280822 245338 280854 245574
rect 280234 209894 280854 245338
rect 280234 209658 280266 209894
rect 280502 209658 280586 209894
rect 280822 209658 280854 209894
rect 280234 209574 280854 209658
rect 280234 209338 280266 209574
rect 280502 209338 280586 209574
rect 280822 209338 280854 209574
rect 280234 173894 280854 209338
rect 280234 173658 280266 173894
rect 280502 173658 280586 173894
rect 280822 173658 280854 173894
rect 280234 173574 280854 173658
rect 280234 173338 280266 173574
rect 280502 173338 280586 173574
rect 280822 173338 280854 173574
rect 280234 137894 280854 173338
rect 280234 137658 280266 137894
rect 280502 137658 280586 137894
rect 280822 137658 280854 137894
rect 280234 137574 280854 137658
rect 280234 137338 280266 137574
rect 280502 137338 280586 137574
rect 280822 137338 280854 137574
rect 280234 101894 280854 137338
rect 280234 101658 280266 101894
rect 280502 101658 280586 101894
rect 280822 101658 280854 101894
rect 280234 101574 280854 101658
rect 280234 101338 280266 101574
rect 280502 101338 280586 101574
rect 280822 101338 280854 101574
rect 280234 65894 280854 101338
rect 280234 65658 280266 65894
rect 280502 65658 280586 65894
rect 280822 65658 280854 65894
rect 280234 65574 280854 65658
rect 280234 65338 280266 65574
rect 280502 65338 280586 65574
rect 280822 65338 280854 65574
rect 280234 29894 280854 65338
rect 280234 29658 280266 29894
rect 280502 29658 280586 29894
rect 280822 29658 280854 29894
rect 280234 29574 280854 29658
rect 280234 29338 280266 29574
rect 280502 29338 280586 29574
rect 280822 29338 280854 29574
rect 280234 -7066 280854 29338
rect 280234 -7302 280266 -7066
rect 280502 -7302 280586 -7066
rect 280822 -7302 280854 -7066
rect 280234 -7386 280854 -7302
rect 280234 -7622 280266 -7386
rect 280502 -7622 280586 -7386
rect 280822 -7622 280854 -7386
rect 280234 -7654 280854 -7622
rect 290194 704838 290814 711590
rect 290194 704602 290226 704838
rect 290462 704602 290546 704838
rect 290782 704602 290814 704838
rect 290194 704518 290814 704602
rect 290194 704282 290226 704518
rect 290462 704282 290546 704518
rect 290782 704282 290814 704518
rect 290194 687854 290814 704282
rect 290194 687618 290226 687854
rect 290462 687618 290546 687854
rect 290782 687618 290814 687854
rect 290194 687534 290814 687618
rect 290194 687298 290226 687534
rect 290462 687298 290546 687534
rect 290782 687298 290814 687534
rect 290194 651854 290814 687298
rect 290194 651618 290226 651854
rect 290462 651618 290546 651854
rect 290782 651618 290814 651854
rect 290194 651534 290814 651618
rect 290194 651298 290226 651534
rect 290462 651298 290546 651534
rect 290782 651298 290814 651534
rect 290194 615854 290814 651298
rect 290194 615618 290226 615854
rect 290462 615618 290546 615854
rect 290782 615618 290814 615854
rect 290194 615534 290814 615618
rect 290194 615298 290226 615534
rect 290462 615298 290546 615534
rect 290782 615298 290814 615534
rect 290194 579854 290814 615298
rect 290194 579618 290226 579854
rect 290462 579618 290546 579854
rect 290782 579618 290814 579854
rect 290194 579534 290814 579618
rect 290194 579298 290226 579534
rect 290462 579298 290546 579534
rect 290782 579298 290814 579534
rect 290194 543854 290814 579298
rect 290194 543618 290226 543854
rect 290462 543618 290546 543854
rect 290782 543618 290814 543854
rect 290194 543534 290814 543618
rect 290194 543298 290226 543534
rect 290462 543298 290546 543534
rect 290782 543298 290814 543534
rect 290194 507854 290814 543298
rect 290194 507618 290226 507854
rect 290462 507618 290546 507854
rect 290782 507618 290814 507854
rect 290194 507534 290814 507618
rect 290194 507298 290226 507534
rect 290462 507298 290546 507534
rect 290782 507298 290814 507534
rect 290194 471854 290814 507298
rect 290194 471618 290226 471854
rect 290462 471618 290546 471854
rect 290782 471618 290814 471854
rect 290194 471534 290814 471618
rect 290194 471298 290226 471534
rect 290462 471298 290546 471534
rect 290782 471298 290814 471534
rect 290194 435854 290814 471298
rect 290194 435618 290226 435854
rect 290462 435618 290546 435854
rect 290782 435618 290814 435854
rect 290194 435534 290814 435618
rect 290194 435298 290226 435534
rect 290462 435298 290546 435534
rect 290782 435298 290814 435534
rect 290194 399854 290814 435298
rect 290194 399618 290226 399854
rect 290462 399618 290546 399854
rect 290782 399618 290814 399854
rect 290194 399534 290814 399618
rect 290194 399298 290226 399534
rect 290462 399298 290546 399534
rect 290782 399298 290814 399534
rect 290194 363854 290814 399298
rect 290194 363618 290226 363854
rect 290462 363618 290546 363854
rect 290782 363618 290814 363854
rect 290194 363534 290814 363618
rect 290194 363298 290226 363534
rect 290462 363298 290546 363534
rect 290782 363298 290814 363534
rect 290194 327854 290814 363298
rect 290194 327618 290226 327854
rect 290462 327618 290546 327854
rect 290782 327618 290814 327854
rect 290194 327534 290814 327618
rect 290194 327298 290226 327534
rect 290462 327298 290546 327534
rect 290782 327298 290814 327534
rect 290194 291854 290814 327298
rect 290194 291618 290226 291854
rect 290462 291618 290546 291854
rect 290782 291618 290814 291854
rect 290194 291534 290814 291618
rect 290194 291298 290226 291534
rect 290462 291298 290546 291534
rect 290782 291298 290814 291534
rect 290194 255854 290814 291298
rect 290194 255618 290226 255854
rect 290462 255618 290546 255854
rect 290782 255618 290814 255854
rect 290194 255534 290814 255618
rect 290194 255298 290226 255534
rect 290462 255298 290546 255534
rect 290782 255298 290814 255534
rect 290194 219854 290814 255298
rect 290194 219618 290226 219854
rect 290462 219618 290546 219854
rect 290782 219618 290814 219854
rect 290194 219534 290814 219618
rect 290194 219298 290226 219534
rect 290462 219298 290546 219534
rect 290782 219298 290814 219534
rect 290194 183854 290814 219298
rect 290194 183618 290226 183854
rect 290462 183618 290546 183854
rect 290782 183618 290814 183854
rect 290194 183534 290814 183618
rect 290194 183298 290226 183534
rect 290462 183298 290546 183534
rect 290782 183298 290814 183534
rect 290194 147854 290814 183298
rect 290194 147618 290226 147854
rect 290462 147618 290546 147854
rect 290782 147618 290814 147854
rect 290194 147534 290814 147618
rect 290194 147298 290226 147534
rect 290462 147298 290546 147534
rect 290782 147298 290814 147534
rect 290194 111854 290814 147298
rect 290194 111618 290226 111854
rect 290462 111618 290546 111854
rect 290782 111618 290814 111854
rect 290194 111534 290814 111618
rect 290194 111298 290226 111534
rect 290462 111298 290546 111534
rect 290782 111298 290814 111534
rect 290194 75854 290814 111298
rect 290194 75618 290226 75854
rect 290462 75618 290546 75854
rect 290782 75618 290814 75854
rect 290194 75534 290814 75618
rect 290194 75298 290226 75534
rect 290462 75298 290546 75534
rect 290782 75298 290814 75534
rect 290194 39854 290814 75298
rect 290194 39618 290226 39854
rect 290462 39618 290546 39854
rect 290782 39618 290814 39854
rect 290194 39534 290814 39618
rect 290194 39298 290226 39534
rect 290462 39298 290546 39534
rect 290782 39298 290814 39534
rect 290194 3854 290814 39298
rect 290194 3618 290226 3854
rect 290462 3618 290546 3854
rect 290782 3618 290814 3854
rect 290194 3534 290814 3618
rect 290194 3298 290226 3534
rect 290462 3298 290546 3534
rect 290782 3298 290814 3534
rect 290194 -346 290814 3298
rect 290194 -582 290226 -346
rect 290462 -582 290546 -346
rect 290782 -582 290814 -346
rect 290194 -666 290814 -582
rect 290194 -902 290226 -666
rect 290462 -902 290546 -666
rect 290782 -902 290814 -666
rect 290194 -7654 290814 -902
rect 293914 705798 294534 711590
rect 293914 705562 293946 705798
rect 294182 705562 294266 705798
rect 294502 705562 294534 705798
rect 293914 705478 294534 705562
rect 293914 705242 293946 705478
rect 294182 705242 294266 705478
rect 294502 705242 294534 705478
rect 293914 691574 294534 705242
rect 293914 691338 293946 691574
rect 294182 691338 294266 691574
rect 294502 691338 294534 691574
rect 293914 691254 294534 691338
rect 293914 691018 293946 691254
rect 294182 691018 294266 691254
rect 294502 691018 294534 691254
rect 293914 655574 294534 691018
rect 293914 655338 293946 655574
rect 294182 655338 294266 655574
rect 294502 655338 294534 655574
rect 293914 655254 294534 655338
rect 293914 655018 293946 655254
rect 294182 655018 294266 655254
rect 294502 655018 294534 655254
rect 293914 619574 294534 655018
rect 293914 619338 293946 619574
rect 294182 619338 294266 619574
rect 294502 619338 294534 619574
rect 293914 619254 294534 619338
rect 293914 619018 293946 619254
rect 294182 619018 294266 619254
rect 294502 619018 294534 619254
rect 293914 583574 294534 619018
rect 293914 583338 293946 583574
rect 294182 583338 294266 583574
rect 294502 583338 294534 583574
rect 293914 583254 294534 583338
rect 293914 583018 293946 583254
rect 294182 583018 294266 583254
rect 294502 583018 294534 583254
rect 293914 547574 294534 583018
rect 293914 547338 293946 547574
rect 294182 547338 294266 547574
rect 294502 547338 294534 547574
rect 293914 547254 294534 547338
rect 293914 547018 293946 547254
rect 294182 547018 294266 547254
rect 294502 547018 294534 547254
rect 293914 511574 294534 547018
rect 293914 511338 293946 511574
rect 294182 511338 294266 511574
rect 294502 511338 294534 511574
rect 293914 511254 294534 511338
rect 293914 511018 293946 511254
rect 294182 511018 294266 511254
rect 294502 511018 294534 511254
rect 293914 475574 294534 511018
rect 293914 475338 293946 475574
rect 294182 475338 294266 475574
rect 294502 475338 294534 475574
rect 293914 475254 294534 475338
rect 293914 475018 293946 475254
rect 294182 475018 294266 475254
rect 294502 475018 294534 475254
rect 293914 439574 294534 475018
rect 293914 439338 293946 439574
rect 294182 439338 294266 439574
rect 294502 439338 294534 439574
rect 293914 439254 294534 439338
rect 293914 439018 293946 439254
rect 294182 439018 294266 439254
rect 294502 439018 294534 439254
rect 293914 403574 294534 439018
rect 293914 403338 293946 403574
rect 294182 403338 294266 403574
rect 294502 403338 294534 403574
rect 293914 403254 294534 403338
rect 293914 403018 293946 403254
rect 294182 403018 294266 403254
rect 294502 403018 294534 403254
rect 293914 367574 294534 403018
rect 293914 367338 293946 367574
rect 294182 367338 294266 367574
rect 294502 367338 294534 367574
rect 293914 367254 294534 367338
rect 293914 367018 293946 367254
rect 294182 367018 294266 367254
rect 294502 367018 294534 367254
rect 293914 331574 294534 367018
rect 293914 331338 293946 331574
rect 294182 331338 294266 331574
rect 294502 331338 294534 331574
rect 293914 331254 294534 331338
rect 293914 331018 293946 331254
rect 294182 331018 294266 331254
rect 294502 331018 294534 331254
rect 293914 295574 294534 331018
rect 293914 295338 293946 295574
rect 294182 295338 294266 295574
rect 294502 295338 294534 295574
rect 293914 295254 294534 295338
rect 293914 295018 293946 295254
rect 294182 295018 294266 295254
rect 294502 295018 294534 295254
rect 293914 259574 294534 295018
rect 293914 259338 293946 259574
rect 294182 259338 294266 259574
rect 294502 259338 294534 259574
rect 293914 259254 294534 259338
rect 293914 259018 293946 259254
rect 294182 259018 294266 259254
rect 294502 259018 294534 259254
rect 293914 223574 294534 259018
rect 293914 223338 293946 223574
rect 294182 223338 294266 223574
rect 294502 223338 294534 223574
rect 293914 223254 294534 223338
rect 293914 223018 293946 223254
rect 294182 223018 294266 223254
rect 294502 223018 294534 223254
rect 293914 187574 294534 223018
rect 293914 187338 293946 187574
rect 294182 187338 294266 187574
rect 294502 187338 294534 187574
rect 293914 187254 294534 187338
rect 293914 187018 293946 187254
rect 294182 187018 294266 187254
rect 294502 187018 294534 187254
rect 293914 151574 294534 187018
rect 293914 151338 293946 151574
rect 294182 151338 294266 151574
rect 294502 151338 294534 151574
rect 293914 151254 294534 151338
rect 293914 151018 293946 151254
rect 294182 151018 294266 151254
rect 294502 151018 294534 151254
rect 293914 115574 294534 151018
rect 293914 115338 293946 115574
rect 294182 115338 294266 115574
rect 294502 115338 294534 115574
rect 293914 115254 294534 115338
rect 293914 115018 293946 115254
rect 294182 115018 294266 115254
rect 294502 115018 294534 115254
rect 293914 79574 294534 115018
rect 293914 79338 293946 79574
rect 294182 79338 294266 79574
rect 294502 79338 294534 79574
rect 293914 79254 294534 79338
rect 293914 79018 293946 79254
rect 294182 79018 294266 79254
rect 294502 79018 294534 79254
rect 293914 43574 294534 79018
rect 293914 43338 293946 43574
rect 294182 43338 294266 43574
rect 294502 43338 294534 43574
rect 293914 43254 294534 43338
rect 293914 43018 293946 43254
rect 294182 43018 294266 43254
rect 294502 43018 294534 43254
rect 293914 7574 294534 43018
rect 297634 706758 298254 711590
rect 297634 706522 297666 706758
rect 297902 706522 297986 706758
rect 298222 706522 298254 706758
rect 297634 706438 298254 706522
rect 297634 706202 297666 706438
rect 297902 706202 297986 706438
rect 298222 706202 298254 706438
rect 297634 695294 298254 706202
rect 297634 695058 297666 695294
rect 297902 695058 297986 695294
rect 298222 695058 298254 695294
rect 297634 694974 298254 695058
rect 297634 694738 297666 694974
rect 297902 694738 297986 694974
rect 298222 694738 298254 694974
rect 297634 659294 298254 694738
rect 297634 659058 297666 659294
rect 297902 659058 297986 659294
rect 298222 659058 298254 659294
rect 297634 658974 298254 659058
rect 297634 658738 297666 658974
rect 297902 658738 297986 658974
rect 298222 658738 298254 658974
rect 297634 623294 298254 658738
rect 297634 623058 297666 623294
rect 297902 623058 297986 623294
rect 298222 623058 298254 623294
rect 297634 622974 298254 623058
rect 297634 622738 297666 622974
rect 297902 622738 297986 622974
rect 298222 622738 298254 622974
rect 297634 587294 298254 622738
rect 297634 587058 297666 587294
rect 297902 587058 297986 587294
rect 298222 587058 298254 587294
rect 297634 586974 298254 587058
rect 297634 586738 297666 586974
rect 297902 586738 297986 586974
rect 298222 586738 298254 586974
rect 297634 551294 298254 586738
rect 297634 551058 297666 551294
rect 297902 551058 297986 551294
rect 298222 551058 298254 551294
rect 297634 550974 298254 551058
rect 297634 550738 297666 550974
rect 297902 550738 297986 550974
rect 298222 550738 298254 550974
rect 297634 515294 298254 550738
rect 297634 515058 297666 515294
rect 297902 515058 297986 515294
rect 298222 515058 298254 515294
rect 297634 514974 298254 515058
rect 297634 514738 297666 514974
rect 297902 514738 297986 514974
rect 298222 514738 298254 514974
rect 297634 479294 298254 514738
rect 297634 479058 297666 479294
rect 297902 479058 297986 479294
rect 298222 479058 298254 479294
rect 297634 478974 298254 479058
rect 297634 478738 297666 478974
rect 297902 478738 297986 478974
rect 298222 478738 298254 478974
rect 297634 443294 298254 478738
rect 297634 443058 297666 443294
rect 297902 443058 297986 443294
rect 298222 443058 298254 443294
rect 297634 442974 298254 443058
rect 297634 442738 297666 442974
rect 297902 442738 297986 442974
rect 298222 442738 298254 442974
rect 297634 407294 298254 442738
rect 297634 407058 297666 407294
rect 297902 407058 297986 407294
rect 298222 407058 298254 407294
rect 297634 406974 298254 407058
rect 297634 406738 297666 406974
rect 297902 406738 297986 406974
rect 298222 406738 298254 406974
rect 297634 371294 298254 406738
rect 297634 371058 297666 371294
rect 297902 371058 297986 371294
rect 298222 371058 298254 371294
rect 297634 370974 298254 371058
rect 297634 370738 297666 370974
rect 297902 370738 297986 370974
rect 298222 370738 298254 370974
rect 297634 335294 298254 370738
rect 297634 335058 297666 335294
rect 297902 335058 297986 335294
rect 298222 335058 298254 335294
rect 297634 334974 298254 335058
rect 297634 334738 297666 334974
rect 297902 334738 297986 334974
rect 298222 334738 298254 334974
rect 297634 299294 298254 334738
rect 297634 299058 297666 299294
rect 297902 299058 297986 299294
rect 298222 299058 298254 299294
rect 297634 298974 298254 299058
rect 297634 298738 297666 298974
rect 297902 298738 297986 298974
rect 298222 298738 298254 298974
rect 297634 263294 298254 298738
rect 297634 263058 297666 263294
rect 297902 263058 297986 263294
rect 298222 263058 298254 263294
rect 297634 262974 298254 263058
rect 297634 262738 297666 262974
rect 297902 262738 297986 262974
rect 298222 262738 298254 262974
rect 297634 227294 298254 262738
rect 297634 227058 297666 227294
rect 297902 227058 297986 227294
rect 298222 227058 298254 227294
rect 297634 226974 298254 227058
rect 297634 226738 297666 226974
rect 297902 226738 297986 226974
rect 298222 226738 298254 226974
rect 297634 191294 298254 226738
rect 297634 191058 297666 191294
rect 297902 191058 297986 191294
rect 298222 191058 298254 191294
rect 297634 190974 298254 191058
rect 297634 190738 297666 190974
rect 297902 190738 297986 190974
rect 298222 190738 298254 190974
rect 297634 155294 298254 190738
rect 297634 155058 297666 155294
rect 297902 155058 297986 155294
rect 298222 155058 298254 155294
rect 297634 154974 298254 155058
rect 297634 154738 297666 154974
rect 297902 154738 297986 154974
rect 298222 154738 298254 154974
rect 297634 119294 298254 154738
rect 297634 119058 297666 119294
rect 297902 119058 297986 119294
rect 298222 119058 298254 119294
rect 297634 118974 298254 119058
rect 297634 118738 297666 118974
rect 297902 118738 297986 118974
rect 298222 118738 298254 118974
rect 297634 83294 298254 118738
rect 297634 83058 297666 83294
rect 297902 83058 297986 83294
rect 298222 83058 298254 83294
rect 297634 82974 298254 83058
rect 297634 82738 297666 82974
rect 297902 82738 297986 82974
rect 298222 82738 298254 82974
rect 297634 47294 298254 82738
rect 297634 47058 297666 47294
rect 297902 47058 297986 47294
rect 298222 47058 298254 47294
rect 297634 46974 298254 47058
rect 297634 46738 297666 46974
rect 297902 46738 297986 46974
rect 298222 46738 298254 46974
rect 297634 11294 298254 46738
rect 297634 11058 297666 11294
rect 297902 11058 297986 11294
rect 298222 11058 298254 11294
rect 297634 10974 298254 11058
rect 297634 10738 297666 10974
rect 297902 10738 297986 10974
rect 298222 10738 298254 10974
rect 293914 7338 293946 7574
rect 294182 7338 294266 7574
rect 294502 7338 294534 7574
rect 293914 7254 294534 7338
rect 293914 7018 293946 7254
rect 294182 7018 294266 7254
rect 294502 7018 294534 7254
rect 293914 -1306 294534 7018
rect 296670 2957 296730 8382
rect 296667 2956 296733 2957
rect 296667 2892 296668 2956
rect 296732 2892 296733 2956
rect 296667 2891 296733 2892
rect 293914 -1542 293946 -1306
rect 294182 -1542 294266 -1306
rect 294502 -1542 294534 -1306
rect 293914 -1626 294534 -1542
rect 293914 -1862 293946 -1626
rect 294182 -1862 294266 -1626
rect 294502 -1862 294534 -1626
rect 293914 -7654 294534 -1862
rect 297634 -2266 298254 10738
rect 297634 -2502 297666 -2266
rect 297902 -2502 297986 -2266
rect 298222 -2502 298254 -2266
rect 297634 -2586 298254 -2502
rect 297634 -2822 297666 -2586
rect 297902 -2822 297986 -2586
rect 298222 -2822 298254 -2586
rect 297634 -7654 298254 -2822
rect 301354 707718 301974 711590
rect 301354 707482 301386 707718
rect 301622 707482 301706 707718
rect 301942 707482 301974 707718
rect 301354 707398 301974 707482
rect 301354 707162 301386 707398
rect 301622 707162 301706 707398
rect 301942 707162 301974 707398
rect 301354 699014 301974 707162
rect 301354 698778 301386 699014
rect 301622 698778 301706 699014
rect 301942 698778 301974 699014
rect 301354 698694 301974 698778
rect 301354 698458 301386 698694
rect 301622 698458 301706 698694
rect 301942 698458 301974 698694
rect 301354 663014 301974 698458
rect 301354 662778 301386 663014
rect 301622 662778 301706 663014
rect 301942 662778 301974 663014
rect 301354 662694 301974 662778
rect 301354 662458 301386 662694
rect 301622 662458 301706 662694
rect 301942 662458 301974 662694
rect 301354 627014 301974 662458
rect 301354 626778 301386 627014
rect 301622 626778 301706 627014
rect 301942 626778 301974 627014
rect 301354 626694 301974 626778
rect 301354 626458 301386 626694
rect 301622 626458 301706 626694
rect 301942 626458 301974 626694
rect 301354 591014 301974 626458
rect 301354 590778 301386 591014
rect 301622 590778 301706 591014
rect 301942 590778 301974 591014
rect 301354 590694 301974 590778
rect 301354 590458 301386 590694
rect 301622 590458 301706 590694
rect 301942 590458 301974 590694
rect 301354 555014 301974 590458
rect 301354 554778 301386 555014
rect 301622 554778 301706 555014
rect 301942 554778 301974 555014
rect 301354 554694 301974 554778
rect 301354 554458 301386 554694
rect 301622 554458 301706 554694
rect 301942 554458 301974 554694
rect 301354 519014 301974 554458
rect 301354 518778 301386 519014
rect 301622 518778 301706 519014
rect 301942 518778 301974 519014
rect 301354 518694 301974 518778
rect 301354 518458 301386 518694
rect 301622 518458 301706 518694
rect 301942 518458 301974 518694
rect 301354 483014 301974 518458
rect 301354 482778 301386 483014
rect 301622 482778 301706 483014
rect 301942 482778 301974 483014
rect 301354 482694 301974 482778
rect 301354 482458 301386 482694
rect 301622 482458 301706 482694
rect 301942 482458 301974 482694
rect 301354 447014 301974 482458
rect 301354 446778 301386 447014
rect 301622 446778 301706 447014
rect 301942 446778 301974 447014
rect 301354 446694 301974 446778
rect 301354 446458 301386 446694
rect 301622 446458 301706 446694
rect 301942 446458 301974 446694
rect 301354 411014 301974 446458
rect 301354 410778 301386 411014
rect 301622 410778 301706 411014
rect 301942 410778 301974 411014
rect 301354 410694 301974 410778
rect 301354 410458 301386 410694
rect 301622 410458 301706 410694
rect 301942 410458 301974 410694
rect 301354 375014 301974 410458
rect 301354 374778 301386 375014
rect 301622 374778 301706 375014
rect 301942 374778 301974 375014
rect 301354 374694 301974 374778
rect 301354 374458 301386 374694
rect 301622 374458 301706 374694
rect 301942 374458 301974 374694
rect 301354 339014 301974 374458
rect 301354 338778 301386 339014
rect 301622 338778 301706 339014
rect 301942 338778 301974 339014
rect 301354 338694 301974 338778
rect 301354 338458 301386 338694
rect 301622 338458 301706 338694
rect 301942 338458 301974 338694
rect 301354 303014 301974 338458
rect 301354 302778 301386 303014
rect 301622 302778 301706 303014
rect 301942 302778 301974 303014
rect 301354 302694 301974 302778
rect 301354 302458 301386 302694
rect 301622 302458 301706 302694
rect 301942 302458 301974 302694
rect 301354 267014 301974 302458
rect 301354 266778 301386 267014
rect 301622 266778 301706 267014
rect 301942 266778 301974 267014
rect 301354 266694 301974 266778
rect 301354 266458 301386 266694
rect 301622 266458 301706 266694
rect 301942 266458 301974 266694
rect 301354 231014 301974 266458
rect 301354 230778 301386 231014
rect 301622 230778 301706 231014
rect 301942 230778 301974 231014
rect 301354 230694 301974 230778
rect 301354 230458 301386 230694
rect 301622 230458 301706 230694
rect 301942 230458 301974 230694
rect 301354 195014 301974 230458
rect 301354 194778 301386 195014
rect 301622 194778 301706 195014
rect 301942 194778 301974 195014
rect 301354 194694 301974 194778
rect 301354 194458 301386 194694
rect 301622 194458 301706 194694
rect 301942 194458 301974 194694
rect 301354 159014 301974 194458
rect 301354 158778 301386 159014
rect 301622 158778 301706 159014
rect 301942 158778 301974 159014
rect 301354 158694 301974 158778
rect 301354 158458 301386 158694
rect 301622 158458 301706 158694
rect 301942 158458 301974 158694
rect 301354 123014 301974 158458
rect 301354 122778 301386 123014
rect 301622 122778 301706 123014
rect 301942 122778 301974 123014
rect 301354 122694 301974 122778
rect 301354 122458 301386 122694
rect 301622 122458 301706 122694
rect 301942 122458 301974 122694
rect 301354 87014 301974 122458
rect 305074 708678 305694 711590
rect 305074 708442 305106 708678
rect 305342 708442 305426 708678
rect 305662 708442 305694 708678
rect 305074 708358 305694 708442
rect 305074 708122 305106 708358
rect 305342 708122 305426 708358
rect 305662 708122 305694 708358
rect 305074 666734 305694 708122
rect 305074 666498 305106 666734
rect 305342 666498 305426 666734
rect 305662 666498 305694 666734
rect 305074 666414 305694 666498
rect 305074 666178 305106 666414
rect 305342 666178 305426 666414
rect 305662 666178 305694 666414
rect 305074 630734 305694 666178
rect 305074 630498 305106 630734
rect 305342 630498 305426 630734
rect 305662 630498 305694 630734
rect 305074 630414 305694 630498
rect 305074 630178 305106 630414
rect 305342 630178 305426 630414
rect 305662 630178 305694 630414
rect 305074 594734 305694 630178
rect 305074 594498 305106 594734
rect 305342 594498 305426 594734
rect 305662 594498 305694 594734
rect 305074 594414 305694 594498
rect 305074 594178 305106 594414
rect 305342 594178 305426 594414
rect 305662 594178 305694 594414
rect 305074 558734 305694 594178
rect 305074 558498 305106 558734
rect 305342 558498 305426 558734
rect 305662 558498 305694 558734
rect 305074 558414 305694 558498
rect 305074 558178 305106 558414
rect 305342 558178 305426 558414
rect 305662 558178 305694 558414
rect 305074 522734 305694 558178
rect 305074 522498 305106 522734
rect 305342 522498 305426 522734
rect 305662 522498 305694 522734
rect 305074 522414 305694 522498
rect 305074 522178 305106 522414
rect 305342 522178 305426 522414
rect 305662 522178 305694 522414
rect 305074 486734 305694 522178
rect 305074 486498 305106 486734
rect 305342 486498 305426 486734
rect 305662 486498 305694 486734
rect 305074 486414 305694 486498
rect 305074 486178 305106 486414
rect 305342 486178 305426 486414
rect 305662 486178 305694 486414
rect 305074 450734 305694 486178
rect 305074 450498 305106 450734
rect 305342 450498 305426 450734
rect 305662 450498 305694 450734
rect 305074 450414 305694 450498
rect 305074 450178 305106 450414
rect 305342 450178 305426 450414
rect 305662 450178 305694 450414
rect 305074 414734 305694 450178
rect 305074 414498 305106 414734
rect 305342 414498 305426 414734
rect 305662 414498 305694 414734
rect 305074 414414 305694 414498
rect 305074 414178 305106 414414
rect 305342 414178 305426 414414
rect 305662 414178 305694 414414
rect 305074 378734 305694 414178
rect 305074 378498 305106 378734
rect 305342 378498 305426 378734
rect 305662 378498 305694 378734
rect 305074 378414 305694 378498
rect 305074 378178 305106 378414
rect 305342 378178 305426 378414
rect 305662 378178 305694 378414
rect 305074 342734 305694 378178
rect 305074 342498 305106 342734
rect 305342 342498 305426 342734
rect 305662 342498 305694 342734
rect 305074 342414 305694 342498
rect 305074 342178 305106 342414
rect 305342 342178 305426 342414
rect 305662 342178 305694 342414
rect 305074 306734 305694 342178
rect 305074 306498 305106 306734
rect 305342 306498 305426 306734
rect 305662 306498 305694 306734
rect 305074 306414 305694 306498
rect 305074 306178 305106 306414
rect 305342 306178 305426 306414
rect 305662 306178 305694 306414
rect 305074 270734 305694 306178
rect 305074 270498 305106 270734
rect 305342 270498 305426 270734
rect 305662 270498 305694 270734
rect 305074 270414 305694 270498
rect 305074 270178 305106 270414
rect 305342 270178 305426 270414
rect 305662 270178 305694 270414
rect 305074 234734 305694 270178
rect 305074 234498 305106 234734
rect 305342 234498 305426 234734
rect 305662 234498 305694 234734
rect 305074 234414 305694 234498
rect 305074 234178 305106 234414
rect 305342 234178 305426 234414
rect 305662 234178 305694 234414
rect 305074 198734 305694 234178
rect 305074 198498 305106 198734
rect 305342 198498 305426 198734
rect 305662 198498 305694 198734
rect 305074 198414 305694 198498
rect 305074 198178 305106 198414
rect 305342 198178 305426 198414
rect 305662 198178 305694 198414
rect 305074 162734 305694 198178
rect 305074 162498 305106 162734
rect 305342 162498 305426 162734
rect 305662 162498 305694 162734
rect 305074 162414 305694 162498
rect 305074 162178 305106 162414
rect 305342 162178 305426 162414
rect 305662 162178 305694 162414
rect 305074 126734 305694 162178
rect 305074 126498 305106 126734
rect 305342 126498 305426 126734
rect 305662 126498 305694 126734
rect 305074 126414 305694 126498
rect 305074 126178 305106 126414
rect 305342 126178 305426 126414
rect 305662 126178 305694 126414
rect 304208 111854 304528 111886
rect 304208 111618 304250 111854
rect 304486 111618 304528 111854
rect 304208 111534 304528 111618
rect 304208 111298 304250 111534
rect 304486 111298 304528 111534
rect 304208 111266 304528 111298
rect 301354 86778 301386 87014
rect 301622 86778 301706 87014
rect 301942 86778 301974 87014
rect 301354 86694 301974 86778
rect 301354 86458 301386 86694
rect 301622 86458 301706 86694
rect 301942 86458 301974 86694
rect 301354 51014 301974 86458
rect 301354 50778 301386 51014
rect 301622 50778 301706 51014
rect 301942 50778 301974 51014
rect 301354 50694 301974 50778
rect 301354 50458 301386 50694
rect 301622 50458 301706 50694
rect 301942 50458 301974 50694
rect 301354 15014 301974 50458
rect 301354 14778 301386 15014
rect 301622 14778 301706 15014
rect 301942 14778 301974 15014
rect 301354 14694 301974 14778
rect 301354 14458 301386 14694
rect 301622 14458 301706 14694
rect 301942 14458 301974 14694
rect 301354 -3226 301974 14458
rect 301354 -3462 301386 -3226
rect 301622 -3462 301706 -3226
rect 301942 -3462 301974 -3226
rect 301354 -3546 301974 -3462
rect 301354 -3782 301386 -3546
rect 301622 -3782 301706 -3546
rect 301942 -3782 301974 -3546
rect 301354 -7654 301974 -3782
rect 305074 90734 305694 126178
rect 305074 90498 305106 90734
rect 305342 90498 305426 90734
rect 305662 90498 305694 90734
rect 305074 90414 305694 90498
rect 305074 90178 305106 90414
rect 305342 90178 305426 90414
rect 305662 90178 305694 90414
rect 305074 54734 305694 90178
rect 305074 54498 305106 54734
rect 305342 54498 305426 54734
rect 305662 54498 305694 54734
rect 305074 54414 305694 54498
rect 305074 54178 305106 54414
rect 305342 54178 305426 54414
rect 305662 54178 305694 54414
rect 305074 18734 305694 54178
rect 305074 18498 305106 18734
rect 305342 18498 305426 18734
rect 305662 18498 305694 18734
rect 305074 18414 305694 18498
rect 305074 18178 305106 18414
rect 305342 18178 305426 18414
rect 305662 18178 305694 18414
rect 305074 -4186 305694 18178
rect 305074 -4422 305106 -4186
rect 305342 -4422 305426 -4186
rect 305662 -4422 305694 -4186
rect 305074 -4506 305694 -4422
rect 305074 -4742 305106 -4506
rect 305342 -4742 305426 -4506
rect 305662 -4742 305694 -4506
rect 305074 -7654 305694 -4742
rect 308794 709638 309414 711590
rect 308794 709402 308826 709638
rect 309062 709402 309146 709638
rect 309382 709402 309414 709638
rect 308794 709318 309414 709402
rect 308794 709082 308826 709318
rect 309062 709082 309146 709318
rect 309382 709082 309414 709318
rect 308794 670454 309414 709082
rect 308794 670218 308826 670454
rect 309062 670218 309146 670454
rect 309382 670218 309414 670454
rect 308794 670134 309414 670218
rect 308794 669898 308826 670134
rect 309062 669898 309146 670134
rect 309382 669898 309414 670134
rect 308794 634454 309414 669898
rect 308794 634218 308826 634454
rect 309062 634218 309146 634454
rect 309382 634218 309414 634454
rect 308794 634134 309414 634218
rect 308794 633898 308826 634134
rect 309062 633898 309146 634134
rect 309382 633898 309414 634134
rect 308794 598454 309414 633898
rect 308794 598218 308826 598454
rect 309062 598218 309146 598454
rect 309382 598218 309414 598454
rect 308794 598134 309414 598218
rect 308794 597898 308826 598134
rect 309062 597898 309146 598134
rect 309382 597898 309414 598134
rect 308794 562454 309414 597898
rect 308794 562218 308826 562454
rect 309062 562218 309146 562454
rect 309382 562218 309414 562454
rect 308794 562134 309414 562218
rect 308794 561898 308826 562134
rect 309062 561898 309146 562134
rect 309382 561898 309414 562134
rect 308794 526454 309414 561898
rect 308794 526218 308826 526454
rect 309062 526218 309146 526454
rect 309382 526218 309414 526454
rect 308794 526134 309414 526218
rect 308794 525898 308826 526134
rect 309062 525898 309146 526134
rect 309382 525898 309414 526134
rect 308794 490454 309414 525898
rect 308794 490218 308826 490454
rect 309062 490218 309146 490454
rect 309382 490218 309414 490454
rect 308794 490134 309414 490218
rect 308794 489898 308826 490134
rect 309062 489898 309146 490134
rect 309382 489898 309414 490134
rect 308794 454454 309414 489898
rect 308794 454218 308826 454454
rect 309062 454218 309146 454454
rect 309382 454218 309414 454454
rect 308794 454134 309414 454218
rect 308794 453898 308826 454134
rect 309062 453898 309146 454134
rect 309382 453898 309414 454134
rect 308794 418454 309414 453898
rect 308794 418218 308826 418454
rect 309062 418218 309146 418454
rect 309382 418218 309414 418454
rect 308794 418134 309414 418218
rect 308794 417898 308826 418134
rect 309062 417898 309146 418134
rect 309382 417898 309414 418134
rect 308794 382454 309414 417898
rect 308794 382218 308826 382454
rect 309062 382218 309146 382454
rect 309382 382218 309414 382454
rect 308794 382134 309414 382218
rect 308794 381898 308826 382134
rect 309062 381898 309146 382134
rect 309382 381898 309414 382134
rect 308794 346454 309414 381898
rect 308794 346218 308826 346454
rect 309062 346218 309146 346454
rect 309382 346218 309414 346454
rect 308794 346134 309414 346218
rect 308794 345898 308826 346134
rect 309062 345898 309146 346134
rect 309382 345898 309414 346134
rect 308794 310454 309414 345898
rect 308794 310218 308826 310454
rect 309062 310218 309146 310454
rect 309382 310218 309414 310454
rect 308794 310134 309414 310218
rect 308794 309898 308826 310134
rect 309062 309898 309146 310134
rect 309382 309898 309414 310134
rect 308794 274454 309414 309898
rect 308794 274218 308826 274454
rect 309062 274218 309146 274454
rect 309382 274218 309414 274454
rect 308794 274134 309414 274218
rect 308794 273898 308826 274134
rect 309062 273898 309146 274134
rect 309382 273898 309414 274134
rect 308794 238454 309414 273898
rect 308794 238218 308826 238454
rect 309062 238218 309146 238454
rect 309382 238218 309414 238454
rect 308794 238134 309414 238218
rect 308794 237898 308826 238134
rect 309062 237898 309146 238134
rect 309382 237898 309414 238134
rect 308794 202454 309414 237898
rect 308794 202218 308826 202454
rect 309062 202218 309146 202454
rect 309382 202218 309414 202454
rect 308794 202134 309414 202218
rect 308794 201898 308826 202134
rect 309062 201898 309146 202134
rect 309382 201898 309414 202134
rect 308794 166454 309414 201898
rect 308794 166218 308826 166454
rect 309062 166218 309146 166454
rect 309382 166218 309414 166454
rect 308794 166134 309414 166218
rect 308794 165898 308826 166134
rect 309062 165898 309146 166134
rect 309382 165898 309414 166134
rect 308794 130454 309414 165898
rect 308794 130218 308826 130454
rect 309062 130218 309146 130454
rect 309382 130218 309414 130454
rect 308794 130134 309414 130218
rect 308794 129898 308826 130134
rect 309062 129898 309146 130134
rect 309382 129898 309414 130134
rect 308794 94454 309414 129898
rect 308794 94218 308826 94454
rect 309062 94218 309146 94454
rect 309382 94218 309414 94454
rect 308794 94134 309414 94218
rect 308794 93898 308826 94134
rect 309062 93898 309146 94134
rect 309382 93898 309414 94134
rect 308794 58454 309414 93898
rect 308794 58218 308826 58454
rect 309062 58218 309146 58454
rect 309382 58218 309414 58454
rect 308794 58134 309414 58218
rect 308794 57898 308826 58134
rect 309062 57898 309146 58134
rect 309382 57898 309414 58134
rect 308794 22454 309414 57898
rect 308794 22218 308826 22454
rect 309062 22218 309146 22454
rect 309382 22218 309414 22454
rect 308794 22134 309414 22218
rect 308794 21898 308826 22134
rect 309062 21898 309146 22134
rect 309382 21898 309414 22134
rect 308794 -5146 309414 21898
rect 308794 -5382 308826 -5146
rect 309062 -5382 309146 -5146
rect 309382 -5382 309414 -5146
rect 308794 -5466 309414 -5382
rect 308794 -5702 308826 -5466
rect 309062 -5702 309146 -5466
rect 309382 -5702 309414 -5466
rect 308794 -7654 309414 -5702
rect 312514 710598 313134 711590
rect 312514 710362 312546 710598
rect 312782 710362 312866 710598
rect 313102 710362 313134 710598
rect 312514 710278 313134 710362
rect 312514 710042 312546 710278
rect 312782 710042 312866 710278
rect 313102 710042 313134 710278
rect 312514 674174 313134 710042
rect 312514 673938 312546 674174
rect 312782 673938 312866 674174
rect 313102 673938 313134 674174
rect 312514 673854 313134 673938
rect 312514 673618 312546 673854
rect 312782 673618 312866 673854
rect 313102 673618 313134 673854
rect 312514 638174 313134 673618
rect 312514 637938 312546 638174
rect 312782 637938 312866 638174
rect 313102 637938 313134 638174
rect 312514 637854 313134 637938
rect 312514 637618 312546 637854
rect 312782 637618 312866 637854
rect 313102 637618 313134 637854
rect 312514 602174 313134 637618
rect 312514 601938 312546 602174
rect 312782 601938 312866 602174
rect 313102 601938 313134 602174
rect 312514 601854 313134 601938
rect 312514 601618 312546 601854
rect 312782 601618 312866 601854
rect 313102 601618 313134 601854
rect 312514 566174 313134 601618
rect 312514 565938 312546 566174
rect 312782 565938 312866 566174
rect 313102 565938 313134 566174
rect 312514 565854 313134 565938
rect 312514 565618 312546 565854
rect 312782 565618 312866 565854
rect 313102 565618 313134 565854
rect 312514 530174 313134 565618
rect 312514 529938 312546 530174
rect 312782 529938 312866 530174
rect 313102 529938 313134 530174
rect 312514 529854 313134 529938
rect 312514 529618 312546 529854
rect 312782 529618 312866 529854
rect 313102 529618 313134 529854
rect 312514 494174 313134 529618
rect 312514 493938 312546 494174
rect 312782 493938 312866 494174
rect 313102 493938 313134 494174
rect 312514 493854 313134 493938
rect 312514 493618 312546 493854
rect 312782 493618 312866 493854
rect 313102 493618 313134 493854
rect 312514 458174 313134 493618
rect 312514 457938 312546 458174
rect 312782 457938 312866 458174
rect 313102 457938 313134 458174
rect 312514 457854 313134 457938
rect 312514 457618 312546 457854
rect 312782 457618 312866 457854
rect 313102 457618 313134 457854
rect 312514 422174 313134 457618
rect 312514 421938 312546 422174
rect 312782 421938 312866 422174
rect 313102 421938 313134 422174
rect 312514 421854 313134 421938
rect 312514 421618 312546 421854
rect 312782 421618 312866 421854
rect 313102 421618 313134 421854
rect 312514 386174 313134 421618
rect 312514 385938 312546 386174
rect 312782 385938 312866 386174
rect 313102 385938 313134 386174
rect 312514 385854 313134 385938
rect 312514 385618 312546 385854
rect 312782 385618 312866 385854
rect 313102 385618 313134 385854
rect 312514 350174 313134 385618
rect 312514 349938 312546 350174
rect 312782 349938 312866 350174
rect 313102 349938 313134 350174
rect 312514 349854 313134 349938
rect 312514 349618 312546 349854
rect 312782 349618 312866 349854
rect 313102 349618 313134 349854
rect 312514 314174 313134 349618
rect 312514 313938 312546 314174
rect 312782 313938 312866 314174
rect 313102 313938 313134 314174
rect 312514 313854 313134 313938
rect 312514 313618 312546 313854
rect 312782 313618 312866 313854
rect 313102 313618 313134 313854
rect 312514 278174 313134 313618
rect 312514 277938 312546 278174
rect 312782 277938 312866 278174
rect 313102 277938 313134 278174
rect 312514 277854 313134 277938
rect 312514 277618 312546 277854
rect 312782 277618 312866 277854
rect 313102 277618 313134 277854
rect 312514 242174 313134 277618
rect 312514 241938 312546 242174
rect 312782 241938 312866 242174
rect 313102 241938 313134 242174
rect 312514 241854 313134 241938
rect 312514 241618 312546 241854
rect 312782 241618 312866 241854
rect 313102 241618 313134 241854
rect 312514 206174 313134 241618
rect 312514 205938 312546 206174
rect 312782 205938 312866 206174
rect 313102 205938 313134 206174
rect 312514 205854 313134 205938
rect 312514 205618 312546 205854
rect 312782 205618 312866 205854
rect 313102 205618 313134 205854
rect 312514 170174 313134 205618
rect 312514 169938 312546 170174
rect 312782 169938 312866 170174
rect 313102 169938 313134 170174
rect 312514 169854 313134 169938
rect 312514 169618 312546 169854
rect 312782 169618 312866 169854
rect 313102 169618 313134 169854
rect 312514 134174 313134 169618
rect 312514 133938 312546 134174
rect 312782 133938 312866 134174
rect 313102 133938 313134 134174
rect 312514 133854 313134 133938
rect 312514 133618 312546 133854
rect 312782 133618 312866 133854
rect 313102 133618 313134 133854
rect 312514 98174 313134 133618
rect 312514 97938 312546 98174
rect 312782 97938 312866 98174
rect 313102 97938 313134 98174
rect 312514 97854 313134 97938
rect 312514 97618 312546 97854
rect 312782 97618 312866 97854
rect 313102 97618 313134 97854
rect 312514 62174 313134 97618
rect 312514 61938 312546 62174
rect 312782 61938 312866 62174
rect 313102 61938 313134 62174
rect 312514 61854 313134 61938
rect 312514 61618 312546 61854
rect 312782 61618 312866 61854
rect 313102 61618 313134 61854
rect 312514 26174 313134 61618
rect 312514 25938 312546 26174
rect 312782 25938 312866 26174
rect 313102 25938 313134 26174
rect 312514 25854 313134 25938
rect 312514 25618 312546 25854
rect 312782 25618 312866 25854
rect 313102 25618 313134 25854
rect 312514 -6106 313134 25618
rect 312514 -6342 312546 -6106
rect 312782 -6342 312866 -6106
rect 313102 -6342 313134 -6106
rect 312514 -6426 313134 -6342
rect 312514 -6662 312546 -6426
rect 312782 -6662 312866 -6426
rect 313102 -6662 313134 -6426
rect 312514 -7654 313134 -6662
rect 316234 711558 316854 711590
rect 316234 711322 316266 711558
rect 316502 711322 316586 711558
rect 316822 711322 316854 711558
rect 316234 711238 316854 711322
rect 316234 711002 316266 711238
rect 316502 711002 316586 711238
rect 316822 711002 316854 711238
rect 316234 677894 316854 711002
rect 316234 677658 316266 677894
rect 316502 677658 316586 677894
rect 316822 677658 316854 677894
rect 316234 677574 316854 677658
rect 316234 677338 316266 677574
rect 316502 677338 316586 677574
rect 316822 677338 316854 677574
rect 316234 641894 316854 677338
rect 316234 641658 316266 641894
rect 316502 641658 316586 641894
rect 316822 641658 316854 641894
rect 316234 641574 316854 641658
rect 316234 641338 316266 641574
rect 316502 641338 316586 641574
rect 316822 641338 316854 641574
rect 316234 605894 316854 641338
rect 316234 605658 316266 605894
rect 316502 605658 316586 605894
rect 316822 605658 316854 605894
rect 316234 605574 316854 605658
rect 316234 605338 316266 605574
rect 316502 605338 316586 605574
rect 316822 605338 316854 605574
rect 316234 569894 316854 605338
rect 316234 569658 316266 569894
rect 316502 569658 316586 569894
rect 316822 569658 316854 569894
rect 316234 569574 316854 569658
rect 316234 569338 316266 569574
rect 316502 569338 316586 569574
rect 316822 569338 316854 569574
rect 316234 533894 316854 569338
rect 316234 533658 316266 533894
rect 316502 533658 316586 533894
rect 316822 533658 316854 533894
rect 316234 533574 316854 533658
rect 316234 533338 316266 533574
rect 316502 533338 316586 533574
rect 316822 533338 316854 533574
rect 316234 497894 316854 533338
rect 316234 497658 316266 497894
rect 316502 497658 316586 497894
rect 316822 497658 316854 497894
rect 316234 497574 316854 497658
rect 316234 497338 316266 497574
rect 316502 497338 316586 497574
rect 316822 497338 316854 497574
rect 316234 461894 316854 497338
rect 316234 461658 316266 461894
rect 316502 461658 316586 461894
rect 316822 461658 316854 461894
rect 316234 461574 316854 461658
rect 316234 461338 316266 461574
rect 316502 461338 316586 461574
rect 316822 461338 316854 461574
rect 316234 425894 316854 461338
rect 316234 425658 316266 425894
rect 316502 425658 316586 425894
rect 316822 425658 316854 425894
rect 316234 425574 316854 425658
rect 316234 425338 316266 425574
rect 316502 425338 316586 425574
rect 316822 425338 316854 425574
rect 316234 389894 316854 425338
rect 316234 389658 316266 389894
rect 316502 389658 316586 389894
rect 316822 389658 316854 389894
rect 316234 389574 316854 389658
rect 316234 389338 316266 389574
rect 316502 389338 316586 389574
rect 316822 389338 316854 389574
rect 316234 353894 316854 389338
rect 316234 353658 316266 353894
rect 316502 353658 316586 353894
rect 316822 353658 316854 353894
rect 316234 353574 316854 353658
rect 316234 353338 316266 353574
rect 316502 353338 316586 353574
rect 316822 353338 316854 353574
rect 316234 317894 316854 353338
rect 316234 317658 316266 317894
rect 316502 317658 316586 317894
rect 316822 317658 316854 317894
rect 316234 317574 316854 317658
rect 316234 317338 316266 317574
rect 316502 317338 316586 317574
rect 316822 317338 316854 317574
rect 316234 281894 316854 317338
rect 316234 281658 316266 281894
rect 316502 281658 316586 281894
rect 316822 281658 316854 281894
rect 316234 281574 316854 281658
rect 316234 281338 316266 281574
rect 316502 281338 316586 281574
rect 316822 281338 316854 281574
rect 316234 245894 316854 281338
rect 316234 245658 316266 245894
rect 316502 245658 316586 245894
rect 316822 245658 316854 245894
rect 316234 245574 316854 245658
rect 316234 245338 316266 245574
rect 316502 245338 316586 245574
rect 316822 245338 316854 245574
rect 316234 209894 316854 245338
rect 316234 209658 316266 209894
rect 316502 209658 316586 209894
rect 316822 209658 316854 209894
rect 316234 209574 316854 209658
rect 316234 209338 316266 209574
rect 316502 209338 316586 209574
rect 316822 209338 316854 209574
rect 316234 173894 316854 209338
rect 316234 173658 316266 173894
rect 316502 173658 316586 173894
rect 316822 173658 316854 173894
rect 316234 173574 316854 173658
rect 316234 173338 316266 173574
rect 316502 173338 316586 173574
rect 316822 173338 316854 173574
rect 316234 137894 316854 173338
rect 316234 137658 316266 137894
rect 316502 137658 316586 137894
rect 316822 137658 316854 137894
rect 316234 137574 316854 137658
rect 316234 137338 316266 137574
rect 316502 137338 316586 137574
rect 316822 137338 316854 137574
rect 316234 101894 316854 137338
rect 326194 704838 326814 711590
rect 326194 704602 326226 704838
rect 326462 704602 326546 704838
rect 326782 704602 326814 704838
rect 326194 704518 326814 704602
rect 326194 704282 326226 704518
rect 326462 704282 326546 704518
rect 326782 704282 326814 704518
rect 326194 687854 326814 704282
rect 326194 687618 326226 687854
rect 326462 687618 326546 687854
rect 326782 687618 326814 687854
rect 326194 687534 326814 687618
rect 326194 687298 326226 687534
rect 326462 687298 326546 687534
rect 326782 687298 326814 687534
rect 326194 651854 326814 687298
rect 326194 651618 326226 651854
rect 326462 651618 326546 651854
rect 326782 651618 326814 651854
rect 326194 651534 326814 651618
rect 326194 651298 326226 651534
rect 326462 651298 326546 651534
rect 326782 651298 326814 651534
rect 326194 615854 326814 651298
rect 326194 615618 326226 615854
rect 326462 615618 326546 615854
rect 326782 615618 326814 615854
rect 326194 615534 326814 615618
rect 326194 615298 326226 615534
rect 326462 615298 326546 615534
rect 326782 615298 326814 615534
rect 326194 579854 326814 615298
rect 326194 579618 326226 579854
rect 326462 579618 326546 579854
rect 326782 579618 326814 579854
rect 326194 579534 326814 579618
rect 326194 579298 326226 579534
rect 326462 579298 326546 579534
rect 326782 579298 326814 579534
rect 326194 543854 326814 579298
rect 326194 543618 326226 543854
rect 326462 543618 326546 543854
rect 326782 543618 326814 543854
rect 326194 543534 326814 543618
rect 326194 543298 326226 543534
rect 326462 543298 326546 543534
rect 326782 543298 326814 543534
rect 326194 507854 326814 543298
rect 326194 507618 326226 507854
rect 326462 507618 326546 507854
rect 326782 507618 326814 507854
rect 326194 507534 326814 507618
rect 326194 507298 326226 507534
rect 326462 507298 326546 507534
rect 326782 507298 326814 507534
rect 326194 471854 326814 507298
rect 326194 471618 326226 471854
rect 326462 471618 326546 471854
rect 326782 471618 326814 471854
rect 326194 471534 326814 471618
rect 326194 471298 326226 471534
rect 326462 471298 326546 471534
rect 326782 471298 326814 471534
rect 326194 435854 326814 471298
rect 326194 435618 326226 435854
rect 326462 435618 326546 435854
rect 326782 435618 326814 435854
rect 326194 435534 326814 435618
rect 326194 435298 326226 435534
rect 326462 435298 326546 435534
rect 326782 435298 326814 435534
rect 326194 399854 326814 435298
rect 326194 399618 326226 399854
rect 326462 399618 326546 399854
rect 326782 399618 326814 399854
rect 326194 399534 326814 399618
rect 326194 399298 326226 399534
rect 326462 399298 326546 399534
rect 326782 399298 326814 399534
rect 326194 363854 326814 399298
rect 326194 363618 326226 363854
rect 326462 363618 326546 363854
rect 326782 363618 326814 363854
rect 326194 363534 326814 363618
rect 326194 363298 326226 363534
rect 326462 363298 326546 363534
rect 326782 363298 326814 363534
rect 326194 327854 326814 363298
rect 326194 327618 326226 327854
rect 326462 327618 326546 327854
rect 326782 327618 326814 327854
rect 326194 327534 326814 327618
rect 326194 327298 326226 327534
rect 326462 327298 326546 327534
rect 326782 327298 326814 327534
rect 326194 291854 326814 327298
rect 326194 291618 326226 291854
rect 326462 291618 326546 291854
rect 326782 291618 326814 291854
rect 326194 291534 326814 291618
rect 326194 291298 326226 291534
rect 326462 291298 326546 291534
rect 326782 291298 326814 291534
rect 326194 255854 326814 291298
rect 326194 255618 326226 255854
rect 326462 255618 326546 255854
rect 326782 255618 326814 255854
rect 326194 255534 326814 255618
rect 326194 255298 326226 255534
rect 326462 255298 326546 255534
rect 326782 255298 326814 255534
rect 326194 219854 326814 255298
rect 326194 219618 326226 219854
rect 326462 219618 326546 219854
rect 326782 219618 326814 219854
rect 326194 219534 326814 219618
rect 326194 219298 326226 219534
rect 326462 219298 326546 219534
rect 326782 219298 326814 219534
rect 326194 183854 326814 219298
rect 326194 183618 326226 183854
rect 326462 183618 326546 183854
rect 326782 183618 326814 183854
rect 326194 183534 326814 183618
rect 326194 183298 326226 183534
rect 326462 183298 326546 183534
rect 326782 183298 326814 183534
rect 326194 147854 326814 183298
rect 326194 147618 326226 147854
rect 326462 147618 326546 147854
rect 326782 147618 326814 147854
rect 326194 147534 326814 147618
rect 326194 147298 326226 147534
rect 326462 147298 326546 147534
rect 326782 147298 326814 147534
rect 319568 115574 319888 115606
rect 319568 115338 319610 115574
rect 319846 115338 319888 115574
rect 319568 115254 319888 115338
rect 319568 115018 319610 115254
rect 319846 115018 319888 115254
rect 319568 114986 319888 115018
rect 316234 101658 316266 101894
rect 316502 101658 316586 101894
rect 316822 101658 316854 101894
rect 316234 101574 316854 101658
rect 316234 101338 316266 101574
rect 316502 101338 316586 101574
rect 316822 101338 316854 101574
rect 316234 65894 316854 101338
rect 326194 111854 326814 147298
rect 326194 111618 326226 111854
rect 326462 111618 326546 111854
rect 326782 111618 326814 111854
rect 326194 111534 326814 111618
rect 326194 111298 326226 111534
rect 326462 111298 326546 111534
rect 326782 111298 326814 111534
rect 324267 78572 324333 78573
rect 324267 78508 324268 78572
rect 324332 78508 324333 78572
rect 324267 78507 324333 78508
rect 324270 77978 324330 78507
rect 316234 65658 316266 65894
rect 316502 65658 316586 65894
rect 316822 65658 316854 65894
rect 316234 65574 316854 65658
rect 316234 65338 316266 65574
rect 316502 65338 316586 65574
rect 316822 65338 316854 65574
rect 316234 29894 316854 65338
rect 316234 29658 316266 29894
rect 316502 29658 316586 29894
rect 316822 29658 316854 29894
rect 316234 29574 316854 29658
rect 316234 29338 316266 29574
rect 316502 29338 316586 29574
rect 316822 29338 316854 29574
rect 316234 -7066 316854 29338
rect 316234 -7302 316266 -7066
rect 316502 -7302 316586 -7066
rect 316822 -7302 316854 -7066
rect 316234 -7386 316854 -7302
rect 316234 -7622 316266 -7386
rect 316502 -7622 316586 -7386
rect 316822 -7622 316854 -7386
rect 316234 -7654 316854 -7622
rect 326194 75854 326814 111298
rect 326194 75618 326226 75854
rect 326462 75618 326546 75854
rect 326782 75618 326814 75854
rect 326194 75534 326814 75618
rect 326194 75298 326226 75534
rect 326462 75298 326546 75534
rect 326782 75298 326814 75534
rect 326194 39854 326814 75298
rect 326194 39618 326226 39854
rect 326462 39618 326546 39854
rect 326782 39618 326814 39854
rect 326194 39534 326814 39618
rect 326194 39298 326226 39534
rect 326462 39298 326546 39534
rect 326782 39298 326814 39534
rect 326194 3854 326814 39298
rect 326194 3618 326226 3854
rect 326462 3618 326546 3854
rect 326782 3618 326814 3854
rect 326194 3534 326814 3618
rect 326194 3298 326226 3534
rect 326462 3298 326546 3534
rect 326782 3298 326814 3534
rect 326194 -346 326814 3298
rect 326194 -582 326226 -346
rect 326462 -582 326546 -346
rect 326782 -582 326814 -346
rect 326194 -666 326814 -582
rect 326194 -902 326226 -666
rect 326462 -902 326546 -666
rect 326782 -902 326814 -666
rect 326194 -7654 326814 -902
rect 329914 705798 330534 711590
rect 329914 705562 329946 705798
rect 330182 705562 330266 705798
rect 330502 705562 330534 705798
rect 329914 705478 330534 705562
rect 329914 705242 329946 705478
rect 330182 705242 330266 705478
rect 330502 705242 330534 705478
rect 329914 691574 330534 705242
rect 329914 691338 329946 691574
rect 330182 691338 330266 691574
rect 330502 691338 330534 691574
rect 329914 691254 330534 691338
rect 329914 691018 329946 691254
rect 330182 691018 330266 691254
rect 330502 691018 330534 691254
rect 329914 655574 330534 691018
rect 329914 655338 329946 655574
rect 330182 655338 330266 655574
rect 330502 655338 330534 655574
rect 329914 655254 330534 655338
rect 329914 655018 329946 655254
rect 330182 655018 330266 655254
rect 330502 655018 330534 655254
rect 329914 619574 330534 655018
rect 329914 619338 329946 619574
rect 330182 619338 330266 619574
rect 330502 619338 330534 619574
rect 329914 619254 330534 619338
rect 329914 619018 329946 619254
rect 330182 619018 330266 619254
rect 330502 619018 330534 619254
rect 329914 583574 330534 619018
rect 329914 583338 329946 583574
rect 330182 583338 330266 583574
rect 330502 583338 330534 583574
rect 329914 583254 330534 583338
rect 329914 583018 329946 583254
rect 330182 583018 330266 583254
rect 330502 583018 330534 583254
rect 329914 547574 330534 583018
rect 329914 547338 329946 547574
rect 330182 547338 330266 547574
rect 330502 547338 330534 547574
rect 329914 547254 330534 547338
rect 329914 547018 329946 547254
rect 330182 547018 330266 547254
rect 330502 547018 330534 547254
rect 329914 511574 330534 547018
rect 329914 511338 329946 511574
rect 330182 511338 330266 511574
rect 330502 511338 330534 511574
rect 329914 511254 330534 511338
rect 329914 511018 329946 511254
rect 330182 511018 330266 511254
rect 330502 511018 330534 511254
rect 329914 475574 330534 511018
rect 329914 475338 329946 475574
rect 330182 475338 330266 475574
rect 330502 475338 330534 475574
rect 329914 475254 330534 475338
rect 329914 475018 329946 475254
rect 330182 475018 330266 475254
rect 330502 475018 330534 475254
rect 329914 439574 330534 475018
rect 329914 439338 329946 439574
rect 330182 439338 330266 439574
rect 330502 439338 330534 439574
rect 329914 439254 330534 439338
rect 329914 439018 329946 439254
rect 330182 439018 330266 439254
rect 330502 439018 330534 439254
rect 329914 403574 330534 439018
rect 329914 403338 329946 403574
rect 330182 403338 330266 403574
rect 330502 403338 330534 403574
rect 329914 403254 330534 403338
rect 329914 403018 329946 403254
rect 330182 403018 330266 403254
rect 330502 403018 330534 403254
rect 329914 367574 330534 403018
rect 329914 367338 329946 367574
rect 330182 367338 330266 367574
rect 330502 367338 330534 367574
rect 329914 367254 330534 367338
rect 329914 367018 329946 367254
rect 330182 367018 330266 367254
rect 330502 367018 330534 367254
rect 329914 331574 330534 367018
rect 329914 331338 329946 331574
rect 330182 331338 330266 331574
rect 330502 331338 330534 331574
rect 329914 331254 330534 331338
rect 329914 331018 329946 331254
rect 330182 331018 330266 331254
rect 330502 331018 330534 331254
rect 329914 295574 330534 331018
rect 329914 295338 329946 295574
rect 330182 295338 330266 295574
rect 330502 295338 330534 295574
rect 329914 295254 330534 295338
rect 329914 295018 329946 295254
rect 330182 295018 330266 295254
rect 330502 295018 330534 295254
rect 329914 259574 330534 295018
rect 329914 259338 329946 259574
rect 330182 259338 330266 259574
rect 330502 259338 330534 259574
rect 329914 259254 330534 259338
rect 329914 259018 329946 259254
rect 330182 259018 330266 259254
rect 330502 259018 330534 259254
rect 329914 223574 330534 259018
rect 329914 223338 329946 223574
rect 330182 223338 330266 223574
rect 330502 223338 330534 223574
rect 329914 223254 330534 223338
rect 329914 223018 329946 223254
rect 330182 223018 330266 223254
rect 330502 223018 330534 223254
rect 329914 187574 330534 223018
rect 329914 187338 329946 187574
rect 330182 187338 330266 187574
rect 330502 187338 330534 187574
rect 329914 187254 330534 187338
rect 329914 187018 329946 187254
rect 330182 187018 330266 187254
rect 330502 187018 330534 187254
rect 329914 151574 330534 187018
rect 329914 151338 329946 151574
rect 330182 151338 330266 151574
rect 330502 151338 330534 151574
rect 329914 151254 330534 151338
rect 329914 151018 329946 151254
rect 330182 151018 330266 151254
rect 330502 151018 330534 151254
rect 329914 115574 330534 151018
rect 329914 115338 329946 115574
rect 330182 115338 330266 115574
rect 330502 115338 330534 115574
rect 329914 115254 330534 115338
rect 329914 115018 329946 115254
rect 330182 115018 330266 115254
rect 330502 115018 330534 115254
rect 329914 79574 330534 115018
rect 329914 79338 329946 79574
rect 330182 79338 330266 79574
rect 330502 79338 330534 79574
rect 329914 79254 330534 79338
rect 329914 79018 329946 79254
rect 330182 79018 330266 79254
rect 330502 79018 330534 79254
rect 329914 43574 330534 79018
rect 329914 43338 329946 43574
rect 330182 43338 330266 43574
rect 330502 43338 330534 43574
rect 329914 43254 330534 43338
rect 329914 43018 329946 43254
rect 330182 43018 330266 43254
rect 330502 43018 330534 43254
rect 329914 7574 330534 43018
rect 329914 7338 329946 7574
rect 330182 7338 330266 7574
rect 330502 7338 330534 7574
rect 329914 7254 330534 7338
rect 329914 7018 329946 7254
rect 330182 7018 330266 7254
rect 330502 7018 330534 7254
rect 329914 -1306 330534 7018
rect 329914 -1542 329946 -1306
rect 330182 -1542 330266 -1306
rect 330502 -1542 330534 -1306
rect 329914 -1626 330534 -1542
rect 329914 -1862 329946 -1626
rect 330182 -1862 330266 -1626
rect 330502 -1862 330534 -1626
rect 329914 -7654 330534 -1862
rect 333634 706758 334254 711590
rect 333634 706522 333666 706758
rect 333902 706522 333986 706758
rect 334222 706522 334254 706758
rect 333634 706438 334254 706522
rect 333634 706202 333666 706438
rect 333902 706202 333986 706438
rect 334222 706202 334254 706438
rect 333634 695294 334254 706202
rect 333634 695058 333666 695294
rect 333902 695058 333986 695294
rect 334222 695058 334254 695294
rect 333634 694974 334254 695058
rect 333634 694738 333666 694974
rect 333902 694738 333986 694974
rect 334222 694738 334254 694974
rect 333634 659294 334254 694738
rect 333634 659058 333666 659294
rect 333902 659058 333986 659294
rect 334222 659058 334254 659294
rect 333634 658974 334254 659058
rect 333634 658738 333666 658974
rect 333902 658738 333986 658974
rect 334222 658738 334254 658974
rect 333634 623294 334254 658738
rect 333634 623058 333666 623294
rect 333902 623058 333986 623294
rect 334222 623058 334254 623294
rect 333634 622974 334254 623058
rect 333634 622738 333666 622974
rect 333902 622738 333986 622974
rect 334222 622738 334254 622974
rect 333634 587294 334254 622738
rect 333634 587058 333666 587294
rect 333902 587058 333986 587294
rect 334222 587058 334254 587294
rect 333634 586974 334254 587058
rect 333634 586738 333666 586974
rect 333902 586738 333986 586974
rect 334222 586738 334254 586974
rect 333634 551294 334254 586738
rect 333634 551058 333666 551294
rect 333902 551058 333986 551294
rect 334222 551058 334254 551294
rect 333634 550974 334254 551058
rect 333634 550738 333666 550974
rect 333902 550738 333986 550974
rect 334222 550738 334254 550974
rect 333634 515294 334254 550738
rect 333634 515058 333666 515294
rect 333902 515058 333986 515294
rect 334222 515058 334254 515294
rect 333634 514974 334254 515058
rect 333634 514738 333666 514974
rect 333902 514738 333986 514974
rect 334222 514738 334254 514974
rect 333634 479294 334254 514738
rect 333634 479058 333666 479294
rect 333902 479058 333986 479294
rect 334222 479058 334254 479294
rect 333634 478974 334254 479058
rect 333634 478738 333666 478974
rect 333902 478738 333986 478974
rect 334222 478738 334254 478974
rect 333634 443294 334254 478738
rect 333634 443058 333666 443294
rect 333902 443058 333986 443294
rect 334222 443058 334254 443294
rect 333634 442974 334254 443058
rect 333634 442738 333666 442974
rect 333902 442738 333986 442974
rect 334222 442738 334254 442974
rect 333634 407294 334254 442738
rect 333634 407058 333666 407294
rect 333902 407058 333986 407294
rect 334222 407058 334254 407294
rect 333634 406974 334254 407058
rect 333634 406738 333666 406974
rect 333902 406738 333986 406974
rect 334222 406738 334254 406974
rect 333634 371294 334254 406738
rect 333634 371058 333666 371294
rect 333902 371058 333986 371294
rect 334222 371058 334254 371294
rect 333634 370974 334254 371058
rect 333634 370738 333666 370974
rect 333902 370738 333986 370974
rect 334222 370738 334254 370974
rect 333634 335294 334254 370738
rect 333634 335058 333666 335294
rect 333902 335058 333986 335294
rect 334222 335058 334254 335294
rect 333634 334974 334254 335058
rect 333634 334738 333666 334974
rect 333902 334738 333986 334974
rect 334222 334738 334254 334974
rect 333634 299294 334254 334738
rect 333634 299058 333666 299294
rect 333902 299058 333986 299294
rect 334222 299058 334254 299294
rect 333634 298974 334254 299058
rect 333634 298738 333666 298974
rect 333902 298738 333986 298974
rect 334222 298738 334254 298974
rect 333634 263294 334254 298738
rect 333634 263058 333666 263294
rect 333902 263058 333986 263294
rect 334222 263058 334254 263294
rect 333634 262974 334254 263058
rect 333634 262738 333666 262974
rect 333902 262738 333986 262974
rect 334222 262738 334254 262974
rect 333634 227294 334254 262738
rect 333634 227058 333666 227294
rect 333902 227058 333986 227294
rect 334222 227058 334254 227294
rect 333634 226974 334254 227058
rect 333634 226738 333666 226974
rect 333902 226738 333986 226974
rect 334222 226738 334254 226974
rect 333634 191294 334254 226738
rect 333634 191058 333666 191294
rect 333902 191058 333986 191294
rect 334222 191058 334254 191294
rect 333634 190974 334254 191058
rect 333634 190738 333666 190974
rect 333902 190738 333986 190974
rect 334222 190738 334254 190974
rect 333634 155294 334254 190738
rect 333634 155058 333666 155294
rect 333902 155058 333986 155294
rect 334222 155058 334254 155294
rect 333634 154974 334254 155058
rect 333634 154738 333666 154974
rect 333902 154738 333986 154974
rect 334222 154738 334254 154974
rect 333634 119294 334254 154738
rect 333634 119058 333666 119294
rect 333902 119058 333986 119294
rect 334222 119058 334254 119294
rect 333634 118974 334254 119058
rect 333634 118738 333666 118974
rect 333902 118738 333986 118974
rect 334222 118738 334254 118974
rect 333634 83294 334254 118738
rect 337354 707718 337974 711590
rect 337354 707482 337386 707718
rect 337622 707482 337706 707718
rect 337942 707482 337974 707718
rect 337354 707398 337974 707482
rect 337354 707162 337386 707398
rect 337622 707162 337706 707398
rect 337942 707162 337974 707398
rect 337354 699014 337974 707162
rect 337354 698778 337386 699014
rect 337622 698778 337706 699014
rect 337942 698778 337974 699014
rect 337354 698694 337974 698778
rect 337354 698458 337386 698694
rect 337622 698458 337706 698694
rect 337942 698458 337974 698694
rect 337354 663014 337974 698458
rect 337354 662778 337386 663014
rect 337622 662778 337706 663014
rect 337942 662778 337974 663014
rect 337354 662694 337974 662778
rect 337354 662458 337386 662694
rect 337622 662458 337706 662694
rect 337942 662458 337974 662694
rect 337354 627014 337974 662458
rect 337354 626778 337386 627014
rect 337622 626778 337706 627014
rect 337942 626778 337974 627014
rect 337354 626694 337974 626778
rect 337354 626458 337386 626694
rect 337622 626458 337706 626694
rect 337942 626458 337974 626694
rect 337354 591014 337974 626458
rect 337354 590778 337386 591014
rect 337622 590778 337706 591014
rect 337942 590778 337974 591014
rect 337354 590694 337974 590778
rect 337354 590458 337386 590694
rect 337622 590458 337706 590694
rect 337942 590458 337974 590694
rect 337354 555014 337974 590458
rect 337354 554778 337386 555014
rect 337622 554778 337706 555014
rect 337942 554778 337974 555014
rect 337354 554694 337974 554778
rect 337354 554458 337386 554694
rect 337622 554458 337706 554694
rect 337942 554458 337974 554694
rect 337354 519014 337974 554458
rect 337354 518778 337386 519014
rect 337622 518778 337706 519014
rect 337942 518778 337974 519014
rect 337354 518694 337974 518778
rect 337354 518458 337386 518694
rect 337622 518458 337706 518694
rect 337942 518458 337974 518694
rect 337354 483014 337974 518458
rect 337354 482778 337386 483014
rect 337622 482778 337706 483014
rect 337942 482778 337974 483014
rect 337354 482694 337974 482778
rect 337354 482458 337386 482694
rect 337622 482458 337706 482694
rect 337942 482458 337974 482694
rect 337354 447014 337974 482458
rect 337354 446778 337386 447014
rect 337622 446778 337706 447014
rect 337942 446778 337974 447014
rect 337354 446694 337974 446778
rect 337354 446458 337386 446694
rect 337622 446458 337706 446694
rect 337942 446458 337974 446694
rect 337354 411014 337974 446458
rect 337354 410778 337386 411014
rect 337622 410778 337706 411014
rect 337942 410778 337974 411014
rect 337354 410694 337974 410778
rect 337354 410458 337386 410694
rect 337622 410458 337706 410694
rect 337942 410458 337974 410694
rect 337354 375014 337974 410458
rect 337354 374778 337386 375014
rect 337622 374778 337706 375014
rect 337942 374778 337974 375014
rect 337354 374694 337974 374778
rect 337354 374458 337386 374694
rect 337622 374458 337706 374694
rect 337942 374458 337974 374694
rect 337354 339014 337974 374458
rect 337354 338778 337386 339014
rect 337622 338778 337706 339014
rect 337942 338778 337974 339014
rect 337354 338694 337974 338778
rect 337354 338458 337386 338694
rect 337622 338458 337706 338694
rect 337942 338458 337974 338694
rect 337354 303014 337974 338458
rect 337354 302778 337386 303014
rect 337622 302778 337706 303014
rect 337942 302778 337974 303014
rect 337354 302694 337974 302778
rect 337354 302458 337386 302694
rect 337622 302458 337706 302694
rect 337942 302458 337974 302694
rect 337354 267014 337974 302458
rect 337354 266778 337386 267014
rect 337622 266778 337706 267014
rect 337942 266778 337974 267014
rect 337354 266694 337974 266778
rect 337354 266458 337386 266694
rect 337622 266458 337706 266694
rect 337942 266458 337974 266694
rect 337354 231014 337974 266458
rect 337354 230778 337386 231014
rect 337622 230778 337706 231014
rect 337942 230778 337974 231014
rect 337354 230694 337974 230778
rect 337354 230458 337386 230694
rect 337622 230458 337706 230694
rect 337942 230458 337974 230694
rect 337354 195014 337974 230458
rect 337354 194778 337386 195014
rect 337622 194778 337706 195014
rect 337942 194778 337974 195014
rect 337354 194694 337974 194778
rect 337354 194458 337386 194694
rect 337622 194458 337706 194694
rect 337942 194458 337974 194694
rect 337354 159014 337974 194458
rect 337354 158778 337386 159014
rect 337622 158778 337706 159014
rect 337942 158778 337974 159014
rect 337354 158694 337974 158778
rect 337354 158458 337386 158694
rect 337622 158458 337706 158694
rect 337942 158458 337974 158694
rect 337354 123014 337974 158458
rect 337354 122778 337386 123014
rect 337622 122778 337706 123014
rect 337942 122778 337974 123014
rect 337354 122694 337974 122778
rect 337354 122458 337386 122694
rect 337622 122458 337706 122694
rect 337942 122458 337974 122694
rect 335859 117468 335925 117469
rect 335859 117404 335860 117468
rect 335924 117404 335925 117468
rect 335859 117403 335925 117404
rect 334928 111854 335248 111886
rect 334928 111618 334970 111854
rect 335206 111618 335248 111854
rect 334928 111534 335248 111618
rect 334928 111298 334970 111534
rect 335206 111298 335248 111534
rect 334928 111266 335248 111298
rect 333634 83058 333666 83294
rect 333902 83058 333986 83294
rect 334222 83058 334254 83294
rect 333634 82974 334254 83058
rect 333634 82738 333666 82974
rect 333902 82738 333986 82974
rect 334222 82738 334254 82974
rect 333634 47294 334254 82738
rect 335675 81292 335741 81293
rect 335675 81228 335676 81292
rect 335740 81228 335741 81292
rect 335675 81227 335741 81228
rect 335678 80613 335738 81227
rect 335675 80612 335741 80613
rect 335675 80548 335676 80612
rect 335740 80548 335741 80612
rect 335675 80547 335741 80548
rect 333634 47058 333666 47294
rect 333902 47058 333986 47294
rect 334222 47058 334254 47294
rect 333634 46974 334254 47058
rect 333634 46738 333666 46974
rect 333902 46738 333986 46974
rect 334222 46738 334254 46974
rect 333634 11294 334254 46738
rect 333634 11058 333666 11294
rect 333902 11058 333986 11294
rect 334222 11058 334254 11294
rect 333634 10974 334254 11058
rect 333634 10738 333666 10974
rect 333902 10738 333986 10974
rect 334222 10738 334254 10974
rect 333634 -2266 334254 10738
rect 335862 8261 335922 117403
rect 336043 116516 336109 116517
rect 336043 116452 336044 116516
rect 336108 116452 336109 116516
rect 336043 116451 336109 116452
rect 336046 8261 336106 116451
rect 336779 110804 336845 110805
rect 336779 110740 336780 110804
rect 336844 110740 336845 110804
rect 336779 110739 336845 110740
rect 336227 107948 336293 107949
rect 336227 107884 336228 107948
rect 336292 107884 336293 107948
rect 336227 107883 336293 107884
rect 335859 8260 335925 8261
rect 335859 8196 335860 8260
rect 335924 8196 335925 8260
rect 335859 8195 335925 8196
rect 336043 8260 336109 8261
rect 336043 8196 336044 8260
rect 336108 8196 336109 8260
rect 336043 8195 336109 8196
rect 336230 8125 336290 107883
rect 336411 98700 336477 98701
rect 336411 98636 336412 98700
rect 336476 98636 336477 98700
rect 336411 98635 336477 98636
rect 336227 8124 336293 8125
rect 336227 8060 336228 8124
rect 336292 8060 336293 8124
rect 336227 8059 336293 8060
rect 336414 7309 336474 98635
rect 336411 7308 336477 7309
rect 336411 7244 336412 7308
rect 336476 7244 336477 7308
rect 336411 7243 336477 7244
rect 336782 6765 336842 110739
rect 337354 87014 337974 122458
rect 341074 708678 341694 711590
rect 341074 708442 341106 708678
rect 341342 708442 341426 708678
rect 341662 708442 341694 708678
rect 341074 708358 341694 708442
rect 341074 708122 341106 708358
rect 341342 708122 341426 708358
rect 341662 708122 341694 708358
rect 341074 666734 341694 708122
rect 341074 666498 341106 666734
rect 341342 666498 341426 666734
rect 341662 666498 341694 666734
rect 341074 666414 341694 666498
rect 341074 666178 341106 666414
rect 341342 666178 341426 666414
rect 341662 666178 341694 666414
rect 341074 630734 341694 666178
rect 341074 630498 341106 630734
rect 341342 630498 341426 630734
rect 341662 630498 341694 630734
rect 341074 630414 341694 630498
rect 341074 630178 341106 630414
rect 341342 630178 341426 630414
rect 341662 630178 341694 630414
rect 341074 594734 341694 630178
rect 341074 594498 341106 594734
rect 341342 594498 341426 594734
rect 341662 594498 341694 594734
rect 341074 594414 341694 594498
rect 341074 594178 341106 594414
rect 341342 594178 341426 594414
rect 341662 594178 341694 594414
rect 341074 558734 341694 594178
rect 341074 558498 341106 558734
rect 341342 558498 341426 558734
rect 341662 558498 341694 558734
rect 341074 558414 341694 558498
rect 341074 558178 341106 558414
rect 341342 558178 341426 558414
rect 341662 558178 341694 558414
rect 341074 522734 341694 558178
rect 341074 522498 341106 522734
rect 341342 522498 341426 522734
rect 341662 522498 341694 522734
rect 341074 522414 341694 522498
rect 341074 522178 341106 522414
rect 341342 522178 341426 522414
rect 341662 522178 341694 522414
rect 341074 486734 341694 522178
rect 341074 486498 341106 486734
rect 341342 486498 341426 486734
rect 341662 486498 341694 486734
rect 341074 486414 341694 486498
rect 341074 486178 341106 486414
rect 341342 486178 341426 486414
rect 341662 486178 341694 486414
rect 341074 450734 341694 486178
rect 341074 450498 341106 450734
rect 341342 450498 341426 450734
rect 341662 450498 341694 450734
rect 341074 450414 341694 450498
rect 341074 450178 341106 450414
rect 341342 450178 341426 450414
rect 341662 450178 341694 450414
rect 341074 414734 341694 450178
rect 341074 414498 341106 414734
rect 341342 414498 341426 414734
rect 341662 414498 341694 414734
rect 341074 414414 341694 414498
rect 341074 414178 341106 414414
rect 341342 414178 341426 414414
rect 341662 414178 341694 414414
rect 341074 378734 341694 414178
rect 341074 378498 341106 378734
rect 341342 378498 341426 378734
rect 341662 378498 341694 378734
rect 341074 378414 341694 378498
rect 341074 378178 341106 378414
rect 341342 378178 341426 378414
rect 341662 378178 341694 378414
rect 341074 342734 341694 378178
rect 341074 342498 341106 342734
rect 341342 342498 341426 342734
rect 341662 342498 341694 342734
rect 341074 342414 341694 342498
rect 341074 342178 341106 342414
rect 341342 342178 341426 342414
rect 341662 342178 341694 342414
rect 341074 306734 341694 342178
rect 341074 306498 341106 306734
rect 341342 306498 341426 306734
rect 341662 306498 341694 306734
rect 341074 306414 341694 306498
rect 341074 306178 341106 306414
rect 341342 306178 341426 306414
rect 341662 306178 341694 306414
rect 341074 270734 341694 306178
rect 341074 270498 341106 270734
rect 341342 270498 341426 270734
rect 341662 270498 341694 270734
rect 341074 270414 341694 270498
rect 341074 270178 341106 270414
rect 341342 270178 341426 270414
rect 341662 270178 341694 270414
rect 341074 234734 341694 270178
rect 341074 234498 341106 234734
rect 341342 234498 341426 234734
rect 341662 234498 341694 234734
rect 341074 234414 341694 234498
rect 341074 234178 341106 234414
rect 341342 234178 341426 234414
rect 341662 234178 341694 234414
rect 341074 198734 341694 234178
rect 341074 198498 341106 198734
rect 341342 198498 341426 198734
rect 341662 198498 341694 198734
rect 341074 198414 341694 198498
rect 341074 198178 341106 198414
rect 341342 198178 341426 198414
rect 341662 198178 341694 198414
rect 341074 162734 341694 198178
rect 341074 162498 341106 162734
rect 341342 162498 341426 162734
rect 341662 162498 341694 162734
rect 341074 162414 341694 162498
rect 341074 162178 341106 162414
rect 341342 162178 341426 162414
rect 341662 162178 341694 162414
rect 341074 126734 341694 162178
rect 341074 126498 341106 126734
rect 341342 126498 341426 126734
rect 341662 126498 341694 126734
rect 341074 126414 341694 126498
rect 341074 126178 341106 126414
rect 341342 126178 341426 126414
rect 341662 126178 341694 126414
rect 338987 111756 339053 111757
rect 338987 111692 338988 111756
rect 339052 111692 339053 111756
rect 338987 111691 339053 111692
rect 338619 109852 338685 109853
rect 338619 109788 338620 109852
rect 338684 109788 338685 109852
rect 338619 109787 338685 109788
rect 338435 106044 338501 106045
rect 338435 105980 338436 106044
rect 338500 105980 338501 106044
rect 338435 105979 338501 105980
rect 337354 86778 337386 87014
rect 337622 86778 337706 87014
rect 337942 86778 337974 87014
rect 337354 86694 337974 86778
rect 337354 86458 337386 86694
rect 337622 86458 337706 86694
rect 337942 86458 337974 86694
rect 337354 51014 337974 86458
rect 337354 50778 337386 51014
rect 337622 50778 337706 51014
rect 337942 50778 337974 51014
rect 337354 50694 337974 50778
rect 337354 50458 337386 50694
rect 337622 50458 337706 50694
rect 337942 50458 337974 50694
rect 337354 15014 337974 50458
rect 337354 14778 337386 15014
rect 337622 14778 337706 15014
rect 337942 14778 337974 15014
rect 337354 14694 337974 14778
rect 337354 14458 337386 14694
rect 337622 14458 337706 14694
rect 337942 14458 337974 14694
rect 336779 6764 336845 6765
rect 336779 6700 336780 6764
rect 336844 6700 336845 6764
rect 336779 6699 336845 6700
rect 335491 3908 335557 3909
rect 335491 3844 335492 3908
rect 335556 3844 335557 3908
rect 335491 3843 335557 3844
rect 335494 3770 335554 3843
rect 335126 3710 335554 3770
rect 335126 3093 335186 3710
rect 335123 3092 335189 3093
rect 335123 3028 335124 3092
rect 335188 3028 335189 3092
rect 335123 3027 335189 3028
rect 333634 -2502 333666 -2266
rect 333902 -2502 333986 -2266
rect 334222 -2502 334254 -2266
rect 333634 -2586 334254 -2502
rect 333634 -2822 333666 -2586
rect 333902 -2822 333986 -2586
rect 334222 -2822 334254 -2586
rect 333634 -7654 334254 -2822
rect 337354 -3226 337974 14458
rect 338438 4538 338498 105979
rect 338622 10437 338682 109787
rect 338803 98428 338869 98429
rect 338803 98364 338804 98428
rect 338868 98364 338869 98428
rect 338803 98363 338869 98364
rect 338619 10436 338685 10437
rect 338619 10372 338620 10436
rect 338684 10372 338685 10436
rect 338619 10371 338685 10372
rect 338806 10301 338866 98363
rect 338803 10300 338869 10301
rect 338803 10236 338804 10300
rect 338868 10236 338869 10300
rect 338803 10235 338869 10236
rect 338990 6578 339050 111691
rect 341074 90734 341694 126178
rect 341074 90498 341106 90734
rect 341342 90498 341426 90734
rect 341662 90498 341694 90734
rect 341074 90414 341694 90498
rect 341074 90178 341106 90414
rect 341342 90178 341426 90414
rect 341662 90178 341694 90414
rect 341074 54734 341694 90178
rect 341074 54498 341106 54734
rect 341342 54498 341426 54734
rect 341662 54498 341694 54734
rect 341074 54414 341694 54498
rect 341074 54178 341106 54414
rect 341342 54178 341426 54414
rect 341662 54178 341694 54414
rect 341074 18734 341694 54178
rect 341074 18498 341106 18734
rect 341342 18498 341426 18734
rect 341662 18498 341694 18734
rect 341074 18414 341694 18498
rect 341074 18178 341106 18414
rect 341342 18178 341426 18414
rect 341662 18178 341694 18414
rect 337354 -3462 337386 -3226
rect 337622 -3462 337706 -3226
rect 337942 -3462 337974 -3226
rect 337354 -3546 337974 -3462
rect 337354 -3782 337386 -3546
rect 337622 -3782 337706 -3546
rect 337942 -3782 337974 -3546
rect 337354 -7654 337974 -3782
rect 341074 -4186 341694 18178
rect 341074 -4422 341106 -4186
rect 341342 -4422 341426 -4186
rect 341662 -4422 341694 -4186
rect 341074 -4506 341694 -4422
rect 341074 -4742 341106 -4506
rect 341342 -4742 341426 -4506
rect 341662 -4742 341694 -4506
rect 341074 -7654 341694 -4742
rect 344794 709638 345414 711590
rect 344794 709402 344826 709638
rect 345062 709402 345146 709638
rect 345382 709402 345414 709638
rect 344794 709318 345414 709402
rect 344794 709082 344826 709318
rect 345062 709082 345146 709318
rect 345382 709082 345414 709318
rect 344794 670454 345414 709082
rect 344794 670218 344826 670454
rect 345062 670218 345146 670454
rect 345382 670218 345414 670454
rect 344794 670134 345414 670218
rect 344794 669898 344826 670134
rect 345062 669898 345146 670134
rect 345382 669898 345414 670134
rect 344794 634454 345414 669898
rect 344794 634218 344826 634454
rect 345062 634218 345146 634454
rect 345382 634218 345414 634454
rect 344794 634134 345414 634218
rect 344794 633898 344826 634134
rect 345062 633898 345146 634134
rect 345382 633898 345414 634134
rect 344794 598454 345414 633898
rect 344794 598218 344826 598454
rect 345062 598218 345146 598454
rect 345382 598218 345414 598454
rect 344794 598134 345414 598218
rect 344794 597898 344826 598134
rect 345062 597898 345146 598134
rect 345382 597898 345414 598134
rect 344794 562454 345414 597898
rect 344794 562218 344826 562454
rect 345062 562218 345146 562454
rect 345382 562218 345414 562454
rect 344794 562134 345414 562218
rect 344794 561898 344826 562134
rect 345062 561898 345146 562134
rect 345382 561898 345414 562134
rect 344794 526454 345414 561898
rect 344794 526218 344826 526454
rect 345062 526218 345146 526454
rect 345382 526218 345414 526454
rect 344794 526134 345414 526218
rect 344794 525898 344826 526134
rect 345062 525898 345146 526134
rect 345382 525898 345414 526134
rect 344794 490454 345414 525898
rect 344794 490218 344826 490454
rect 345062 490218 345146 490454
rect 345382 490218 345414 490454
rect 344794 490134 345414 490218
rect 344794 489898 344826 490134
rect 345062 489898 345146 490134
rect 345382 489898 345414 490134
rect 344794 454454 345414 489898
rect 344794 454218 344826 454454
rect 345062 454218 345146 454454
rect 345382 454218 345414 454454
rect 344794 454134 345414 454218
rect 344794 453898 344826 454134
rect 345062 453898 345146 454134
rect 345382 453898 345414 454134
rect 344794 418454 345414 453898
rect 344794 418218 344826 418454
rect 345062 418218 345146 418454
rect 345382 418218 345414 418454
rect 344794 418134 345414 418218
rect 344794 417898 344826 418134
rect 345062 417898 345146 418134
rect 345382 417898 345414 418134
rect 344794 382454 345414 417898
rect 344794 382218 344826 382454
rect 345062 382218 345146 382454
rect 345382 382218 345414 382454
rect 344794 382134 345414 382218
rect 344794 381898 344826 382134
rect 345062 381898 345146 382134
rect 345382 381898 345414 382134
rect 344794 346454 345414 381898
rect 344794 346218 344826 346454
rect 345062 346218 345146 346454
rect 345382 346218 345414 346454
rect 344794 346134 345414 346218
rect 344794 345898 344826 346134
rect 345062 345898 345146 346134
rect 345382 345898 345414 346134
rect 344794 310454 345414 345898
rect 344794 310218 344826 310454
rect 345062 310218 345146 310454
rect 345382 310218 345414 310454
rect 344794 310134 345414 310218
rect 344794 309898 344826 310134
rect 345062 309898 345146 310134
rect 345382 309898 345414 310134
rect 344794 274454 345414 309898
rect 344794 274218 344826 274454
rect 345062 274218 345146 274454
rect 345382 274218 345414 274454
rect 344794 274134 345414 274218
rect 344794 273898 344826 274134
rect 345062 273898 345146 274134
rect 345382 273898 345414 274134
rect 344794 238454 345414 273898
rect 344794 238218 344826 238454
rect 345062 238218 345146 238454
rect 345382 238218 345414 238454
rect 344794 238134 345414 238218
rect 344794 237898 344826 238134
rect 345062 237898 345146 238134
rect 345382 237898 345414 238134
rect 344794 202454 345414 237898
rect 344794 202218 344826 202454
rect 345062 202218 345146 202454
rect 345382 202218 345414 202454
rect 344794 202134 345414 202218
rect 344794 201898 344826 202134
rect 345062 201898 345146 202134
rect 345382 201898 345414 202134
rect 344794 166454 345414 201898
rect 344794 166218 344826 166454
rect 345062 166218 345146 166454
rect 345382 166218 345414 166454
rect 344794 166134 345414 166218
rect 344794 165898 344826 166134
rect 345062 165898 345146 166134
rect 345382 165898 345414 166134
rect 344794 130454 345414 165898
rect 344794 130218 344826 130454
rect 345062 130218 345146 130454
rect 345382 130218 345414 130454
rect 344794 130134 345414 130218
rect 344794 129898 344826 130134
rect 345062 129898 345146 130134
rect 345382 129898 345414 130134
rect 344794 94454 345414 129898
rect 344794 94218 344826 94454
rect 345062 94218 345146 94454
rect 345382 94218 345414 94454
rect 344794 94134 345414 94218
rect 344794 93898 344826 94134
rect 345062 93898 345146 94134
rect 345382 93898 345414 94134
rect 344794 58454 345414 93898
rect 344794 58218 344826 58454
rect 345062 58218 345146 58454
rect 345382 58218 345414 58454
rect 344794 58134 345414 58218
rect 344794 57898 344826 58134
rect 345062 57898 345146 58134
rect 345382 57898 345414 58134
rect 344794 22454 345414 57898
rect 344794 22218 344826 22454
rect 345062 22218 345146 22454
rect 345382 22218 345414 22454
rect 344794 22134 345414 22218
rect 344794 21898 344826 22134
rect 345062 21898 345146 22134
rect 345382 21898 345414 22134
rect 344794 -5146 345414 21898
rect 344794 -5382 344826 -5146
rect 345062 -5382 345146 -5146
rect 345382 -5382 345414 -5146
rect 344794 -5466 345414 -5382
rect 344794 -5702 344826 -5466
rect 345062 -5702 345146 -5466
rect 345382 -5702 345414 -5466
rect 344794 -7654 345414 -5702
rect 348514 710598 349134 711590
rect 348514 710362 348546 710598
rect 348782 710362 348866 710598
rect 349102 710362 349134 710598
rect 348514 710278 349134 710362
rect 348514 710042 348546 710278
rect 348782 710042 348866 710278
rect 349102 710042 349134 710278
rect 348514 674174 349134 710042
rect 348514 673938 348546 674174
rect 348782 673938 348866 674174
rect 349102 673938 349134 674174
rect 348514 673854 349134 673938
rect 348514 673618 348546 673854
rect 348782 673618 348866 673854
rect 349102 673618 349134 673854
rect 348514 638174 349134 673618
rect 348514 637938 348546 638174
rect 348782 637938 348866 638174
rect 349102 637938 349134 638174
rect 348514 637854 349134 637938
rect 348514 637618 348546 637854
rect 348782 637618 348866 637854
rect 349102 637618 349134 637854
rect 348514 602174 349134 637618
rect 348514 601938 348546 602174
rect 348782 601938 348866 602174
rect 349102 601938 349134 602174
rect 348514 601854 349134 601938
rect 348514 601618 348546 601854
rect 348782 601618 348866 601854
rect 349102 601618 349134 601854
rect 348514 566174 349134 601618
rect 348514 565938 348546 566174
rect 348782 565938 348866 566174
rect 349102 565938 349134 566174
rect 348514 565854 349134 565938
rect 348514 565618 348546 565854
rect 348782 565618 348866 565854
rect 349102 565618 349134 565854
rect 348514 530174 349134 565618
rect 348514 529938 348546 530174
rect 348782 529938 348866 530174
rect 349102 529938 349134 530174
rect 348514 529854 349134 529938
rect 348514 529618 348546 529854
rect 348782 529618 348866 529854
rect 349102 529618 349134 529854
rect 348514 494174 349134 529618
rect 348514 493938 348546 494174
rect 348782 493938 348866 494174
rect 349102 493938 349134 494174
rect 348514 493854 349134 493938
rect 348514 493618 348546 493854
rect 348782 493618 348866 493854
rect 349102 493618 349134 493854
rect 348514 458174 349134 493618
rect 348514 457938 348546 458174
rect 348782 457938 348866 458174
rect 349102 457938 349134 458174
rect 348514 457854 349134 457938
rect 348514 457618 348546 457854
rect 348782 457618 348866 457854
rect 349102 457618 349134 457854
rect 348514 422174 349134 457618
rect 348514 421938 348546 422174
rect 348782 421938 348866 422174
rect 349102 421938 349134 422174
rect 348514 421854 349134 421938
rect 348514 421618 348546 421854
rect 348782 421618 348866 421854
rect 349102 421618 349134 421854
rect 348514 386174 349134 421618
rect 348514 385938 348546 386174
rect 348782 385938 348866 386174
rect 349102 385938 349134 386174
rect 348514 385854 349134 385938
rect 348514 385618 348546 385854
rect 348782 385618 348866 385854
rect 349102 385618 349134 385854
rect 348514 350174 349134 385618
rect 348514 349938 348546 350174
rect 348782 349938 348866 350174
rect 349102 349938 349134 350174
rect 348514 349854 349134 349938
rect 348514 349618 348546 349854
rect 348782 349618 348866 349854
rect 349102 349618 349134 349854
rect 348514 314174 349134 349618
rect 348514 313938 348546 314174
rect 348782 313938 348866 314174
rect 349102 313938 349134 314174
rect 348514 313854 349134 313938
rect 348514 313618 348546 313854
rect 348782 313618 348866 313854
rect 349102 313618 349134 313854
rect 348514 278174 349134 313618
rect 348514 277938 348546 278174
rect 348782 277938 348866 278174
rect 349102 277938 349134 278174
rect 348514 277854 349134 277938
rect 348514 277618 348546 277854
rect 348782 277618 348866 277854
rect 349102 277618 349134 277854
rect 348514 242174 349134 277618
rect 348514 241938 348546 242174
rect 348782 241938 348866 242174
rect 349102 241938 349134 242174
rect 348514 241854 349134 241938
rect 348514 241618 348546 241854
rect 348782 241618 348866 241854
rect 349102 241618 349134 241854
rect 348514 206174 349134 241618
rect 348514 205938 348546 206174
rect 348782 205938 348866 206174
rect 349102 205938 349134 206174
rect 348514 205854 349134 205938
rect 348514 205618 348546 205854
rect 348782 205618 348866 205854
rect 349102 205618 349134 205854
rect 348514 170174 349134 205618
rect 348514 169938 348546 170174
rect 348782 169938 348866 170174
rect 349102 169938 349134 170174
rect 348514 169854 349134 169938
rect 348514 169618 348546 169854
rect 348782 169618 348866 169854
rect 349102 169618 349134 169854
rect 348514 134174 349134 169618
rect 348514 133938 348546 134174
rect 348782 133938 348866 134174
rect 349102 133938 349134 134174
rect 348514 133854 349134 133938
rect 348514 133618 348546 133854
rect 348782 133618 348866 133854
rect 349102 133618 349134 133854
rect 348514 98174 349134 133618
rect 348514 97938 348546 98174
rect 348782 97938 348866 98174
rect 349102 97938 349134 98174
rect 348514 97854 349134 97938
rect 348514 97618 348546 97854
rect 348782 97618 348866 97854
rect 349102 97618 349134 97854
rect 348514 62174 349134 97618
rect 348514 61938 348546 62174
rect 348782 61938 348866 62174
rect 349102 61938 349134 62174
rect 348514 61854 349134 61938
rect 348514 61618 348546 61854
rect 348782 61618 348866 61854
rect 349102 61618 349134 61854
rect 348514 26174 349134 61618
rect 348514 25938 348546 26174
rect 348782 25938 348866 26174
rect 349102 25938 349134 26174
rect 348514 25854 349134 25938
rect 348514 25618 348546 25854
rect 348782 25618 348866 25854
rect 349102 25618 349134 25854
rect 348514 -6106 349134 25618
rect 348514 -6342 348546 -6106
rect 348782 -6342 348866 -6106
rect 349102 -6342 349134 -6106
rect 348514 -6426 349134 -6342
rect 348514 -6662 348546 -6426
rect 348782 -6662 348866 -6426
rect 349102 -6662 349134 -6426
rect 348514 -7654 349134 -6662
rect 352234 711558 352854 711590
rect 352234 711322 352266 711558
rect 352502 711322 352586 711558
rect 352822 711322 352854 711558
rect 352234 711238 352854 711322
rect 352234 711002 352266 711238
rect 352502 711002 352586 711238
rect 352822 711002 352854 711238
rect 352234 677894 352854 711002
rect 352234 677658 352266 677894
rect 352502 677658 352586 677894
rect 352822 677658 352854 677894
rect 352234 677574 352854 677658
rect 352234 677338 352266 677574
rect 352502 677338 352586 677574
rect 352822 677338 352854 677574
rect 352234 641894 352854 677338
rect 352234 641658 352266 641894
rect 352502 641658 352586 641894
rect 352822 641658 352854 641894
rect 352234 641574 352854 641658
rect 352234 641338 352266 641574
rect 352502 641338 352586 641574
rect 352822 641338 352854 641574
rect 352234 605894 352854 641338
rect 352234 605658 352266 605894
rect 352502 605658 352586 605894
rect 352822 605658 352854 605894
rect 352234 605574 352854 605658
rect 352234 605338 352266 605574
rect 352502 605338 352586 605574
rect 352822 605338 352854 605574
rect 352234 569894 352854 605338
rect 352234 569658 352266 569894
rect 352502 569658 352586 569894
rect 352822 569658 352854 569894
rect 352234 569574 352854 569658
rect 352234 569338 352266 569574
rect 352502 569338 352586 569574
rect 352822 569338 352854 569574
rect 352234 533894 352854 569338
rect 352234 533658 352266 533894
rect 352502 533658 352586 533894
rect 352822 533658 352854 533894
rect 352234 533574 352854 533658
rect 352234 533338 352266 533574
rect 352502 533338 352586 533574
rect 352822 533338 352854 533574
rect 352234 497894 352854 533338
rect 352234 497658 352266 497894
rect 352502 497658 352586 497894
rect 352822 497658 352854 497894
rect 352234 497574 352854 497658
rect 352234 497338 352266 497574
rect 352502 497338 352586 497574
rect 352822 497338 352854 497574
rect 352234 461894 352854 497338
rect 352234 461658 352266 461894
rect 352502 461658 352586 461894
rect 352822 461658 352854 461894
rect 352234 461574 352854 461658
rect 352234 461338 352266 461574
rect 352502 461338 352586 461574
rect 352822 461338 352854 461574
rect 352234 425894 352854 461338
rect 352234 425658 352266 425894
rect 352502 425658 352586 425894
rect 352822 425658 352854 425894
rect 352234 425574 352854 425658
rect 352234 425338 352266 425574
rect 352502 425338 352586 425574
rect 352822 425338 352854 425574
rect 352234 389894 352854 425338
rect 352234 389658 352266 389894
rect 352502 389658 352586 389894
rect 352822 389658 352854 389894
rect 352234 389574 352854 389658
rect 352234 389338 352266 389574
rect 352502 389338 352586 389574
rect 352822 389338 352854 389574
rect 352234 353894 352854 389338
rect 352234 353658 352266 353894
rect 352502 353658 352586 353894
rect 352822 353658 352854 353894
rect 352234 353574 352854 353658
rect 352234 353338 352266 353574
rect 352502 353338 352586 353574
rect 352822 353338 352854 353574
rect 352234 317894 352854 353338
rect 352234 317658 352266 317894
rect 352502 317658 352586 317894
rect 352822 317658 352854 317894
rect 352234 317574 352854 317658
rect 352234 317338 352266 317574
rect 352502 317338 352586 317574
rect 352822 317338 352854 317574
rect 352234 281894 352854 317338
rect 352234 281658 352266 281894
rect 352502 281658 352586 281894
rect 352822 281658 352854 281894
rect 352234 281574 352854 281658
rect 352234 281338 352266 281574
rect 352502 281338 352586 281574
rect 352822 281338 352854 281574
rect 352234 245894 352854 281338
rect 352234 245658 352266 245894
rect 352502 245658 352586 245894
rect 352822 245658 352854 245894
rect 352234 245574 352854 245658
rect 352234 245338 352266 245574
rect 352502 245338 352586 245574
rect 352822 245338 352854 245574
rect 352234 209894 352854 245338
rect 352234 209658 352266 209894
rect 352502 209658 352586 209894
rect 352822 209658 352854 209894
rect 352234 209574 352854 209658
rect 352234 209338 352266 209574
rect 352502 209338 352586 209574
rect 352822 209338 352854 209574
rect 352234 173894 352854 209338
rect 352234 173658 352266 173894
rect 352502 173658 352586 173894
rect 352822 173658 352854 173894
rect 352234 173574 352854 173658
rect 352234 173338 352266 173574
rect 352502 173338 352586 173574
rect 352822 173338 352854 173574
rect 352234 137894 352854 173338
rect 352234 137658 352266 137894
rect 352502 137658 352586 137894
rect 352822 137658 352854 137894
rect 352234 137574 352854 137658
rect 352234 137338 352266 137574
rect 352502 137338 352586 137574
rect 352822 137338 352854 137574
rect 352234 101894 352854 137338
rect 352234 101658 352266 101894
rect 352502 101658 352586 101894
rect 352822 101658 352854 101894
rect 352234 101574 352854 101658
rect 352234 101338 352266 101574
rect 352502 101338 352586 101574
rect 352822 101338 352854 101574
rect 352234 65894 352854 101338
rect 352234 65658 352266 65894
rect 352502 65658 352586 65894
rect 352822 65658 352854 65894
rect 352234 65574 352854 65658
rect 352234 65338 352266 65574
rect 352502 65338 352586 65574
rect 352822 65338 352854 65574
rect 352234 29894 352854 65338
rect 352234 29658 352266 29894
rect 352502 29658 352586 29894
rect 352822 29658 352854 29894
rect 352234 29574 352854 29658
rect 352234 29338 352266 29574
rect 352502 29338 352586 29574
rect 352822 29338 352854 29574
rect 352234 -7066 352854 29338
rect 352234 -7302 352266 -7066
rect 352502 -7302 352586 -7066
rect 352822 -7302 352854 -7066
rect 352234 -7386 352854 -7302
rect 352234 -7622 352266 -7386
rect 352502 -7622 352586 -7386
rect 352822 -7622 352854 -7386
rect 352234 -7654 352854 -7622
rect 362194 704838 362814 711590
rect 362194 704602 362226 704838
rect 362462 704602 362546 704838
rect 362782 704602 362814 704838
rect 362194 704518 362814 704602
rect 362194 704282 362226 704518
rect 362462 704282 362546 704518
rect 362782 704282 362814 704518
rect 362194 687854 362814 704282
rect 362194 687618 362226 687854
rect 362462 687618 362546 687854
rect 362782 687618 362814 687854
rect 362194 687534 362814 687618
rect 362194 687298 362226 687534
rect 362462 687298 362546 687534
rect 362782 687298 362814 687534
rect 362194 651854 362814 687298
rect 362194 651618 362226 651854
rect 362462 651618 362546 651854
rect 362782 651618 362814 651854
rect 362194 651534 362814 651618
rect 362194 651298 362226 651534
rect 362462 651298 362546 651534
rect 362782 651298 362814 651534
rect 362194 615854 362814 651298
rect 362194 615618 362226 615854
rect 362462 615618 362546 615854
rect 362782 615618 362814 615854
rect 362194 615534 362814 615618
rect 362194 615298 362226 615534
rect 362462 615298 362546 615534
rect 362782 615298 362814 615534
rect 362194 579854 362814 615298
rect 362194 579618 362226 579854
rect 362462 579618 362546 579854
rect 362782 579618 362814 579854
rect 362194 579534 362814 579618
rect 362194 579298 362226 579534
rect 362462 579298 362546 579534
rect 362782 579298 362814 579534
rect 362194 543854 362814 579298
rect 362194 543618 362226 543854
rect 362462 543618 362546 543854
rect 362782 543618 362814 543854
rect 362194 543534 362814 543618
rect 362194 543298 362226 543534
rect 362462 543298 362546 543534
rect 362782 543298 362814 543534
rect 362194 507854 362814 543298
rect 362194 507618 362226 507854
rect 362462 507618 362546 507854
rect 362782 507618 362814 507854
rect 362194 507534 362814 507618
rect 362194 507298 362226 507534
rect 362462 507298 362546 507534
rect 362782 507298 362814 507534
rect 362194 471854 362814 507298
rect 362194 471618 362226 471854
rect 362462 471618 362546 471854
rect 362782 471618 362814 471854
rect 362194 471534 362814 471618
rect 362194 471298 362226 471534
rect 362462 471298 362546 471534
rect 362782 471298 362814 471534
rect 362194 435854 362814 471298
rect 362194 435618 362226 435854
rect 362462 435618 362546 435854
rect 362782 435618 362814 435854
rect 362194 435534 362814 435618
rect 362194 435298 362226 435534
rect 362462 435298 362546 435534
rect 362782 435298 362814 435534
rect 362194 399854 362814 435298
rect 362194 399618 362226 399854
rect 362462 399618 362546 399854
rect 362782 399618 362814 399854
rect 362194 399534 362814 399618
rect 362194 399298 362226 399534
rect 362462 399298 362546 399534
rect 362782 399298 362814 399534
rect 362194 363854 362814 399298
rect 362194 363618 362226 363854
rect 362462 363618 362546 363854
rect 362782 363618 362814 363854
rect 362194 363534 362814 363618
rect 362194 363298 362226 363534
rect 362462 363298 362546 363534
rect 362782 363298 362814 363534
rect 362194 327854 362814 363298
rect 362194 327618 362226 327854
rect 362462 327618 362546 327854
rect 362782 327618 362814 327854
rect 362194 327534 362814 327618
rect 362194 327298 362226 327534
rect 362462 327298 362546 327534
rect 362782 327298 362814 327534
rect 362194 291854 362814 327298
rect 362194 291618 362226 291854
rect 362462 291618 362546 291854
rect 362782 291618 362814 291854
rect 362194 291534 362814 291618
rect 362194 291298 362226 291534
rect 362462 291298 362546 291534
rect 362782 291298 362814 291534
rect 362194 255854 362814 291298
rect 362194 255618 362226 255854
rect 362462 255618 362546 255854
rect 362782 255618 362814 255854
rect 362194 255534 362814 255618
rect 362194 255298 362226 255534
rect 362462 255298 362546 255534
rect 362782 255298 362814 255534
rect 362194 219854 362814 255298
rect 362194 219618 362226 219854
rect 362462 219618 362546 219854
rect 362782 219618 362814 219854
rect 362194 219534 362814 219618
rect 362194 219298 362226 219534
rect 362462 219298 362546 219534
rect 362782 219298 362814 219534
rect 362194 183854 362814 219298
rect 362194 183618 362226 183854
rect 362462 183618 362546 183854
rect 362782 183618 362814 183854
rect 362194 183534 362814 183618
rect 362194 183298 362226 183534
rect 362462 183298 362546 183534
rect 362782 183298 362814 183534
rect 362194 147854 362814 183298
rect 362194 147618 362226 147854
rect 362462 147618 362546 147854
rect 362782 147618 362814 147854
rect 362194 147534 362814 147618
rect 362194 147298 362226 147534
rect 362462 147298 362546 147534
rect 362782 147298 362814 147534
rect 362194 111854 362814 147298
rect 362194 111618 362226 111854
rect 362462 111618 362546 111854
rect 362782 111618 362814 111854
rect 362194 111534 362814 111618
rect 362194 111298 362226 111534
rect 362462 111298 362546 111534
rect 362782 111298 362814 111534
rect 362194 75854 362814 111298
rect 362194 75618 362226 75854
rect 362462 75618 362546 75854
rect 362782 75618 362814 75854
rect 362194 75534 362814 75618
rect 362194 75298 362226 75534
rect 362462 75298 362546 75534
rect 362782 75298 362814 75534
rect 362194 39854 362814 75298
rect 362194 39618 362226 39854
rect 362462 39618 362546 39854
rect 362782 39618 362814 39854
rect 362194 39534 362814 39618
rect 362194 39298 362226 39534
rect 362462 39298 362546 39534
rect 362782 39298 362814 39534
rect 362194 3854 362814 39298
rect 362194 3618 362226 3854
rect 362462 3618 362546 3854
rect 362782 3618 362814 3854
rect 362194 3534 362814 3618
rect 362194 3298 362226 3534
rect 362462 3298 362546 3534
rect 362782 3298 362814 3534
rect 362194 -346 362814 3298
rect 362194 -582 362226 -346
rect 362462 -582 362546 -346
rect 362782 -582 362814 -346
rect 362194 -666 362814 -582
rect 362194 -902 362226 -666
rect 362462 -902 362546 -666
rect 362782 -902 362814 -666
rect 362194 -7654 362814 -902
rect 365914 705798 366534 711590
rect 365914 705562 365946 705798
rect 366182 705562 366266 705798
rect 366502 705562 366534 705798
rect 365914 705478 366534 705562
rect 365914 705242 365946 705478
rect 366182 705242 366266 705478
rect 366502 705242 366534 705478
rect 365914 691574 366534 705242
rect 365914 691338 365946 691574
rect 366182 691338 366266 691574
rect 366502 691338 366534 691574
rect 365914 691254 366534 691338
rect 365914 691018 365946 691254
rect 366182 691018 366266 691254
rect 366502 691018 366534 691254
rect 365914 655574 366534 691018
rect 365914 655338 365946 655574
rect 366182 655338 366266 655574
rect 366502 655338 366534 655574
rect 365914 655254 366534 655338
rect 365914 655018 365946 655254
rect 366182 655018 366266 655254
rect 366502 655018 366534 655254
rect 365914 619574 366534 655018
rect 365914 619338 365946 619574
rect 366182 619338 366266 619574
rect 366502 619338 366534 619574
rect 365914 619254 366534 619338
rect 365914 619018 365946 619254
rect 366182 619018 366266 619254
rect 366502 619018 366534 619254
rect 365914 583574 366534 619018
rect 365914 583338 365946 583574
rect 366182 583338 366266 583574
rect 366502 583338 366534 583574
rect 365914 583254 366534 583338
rect 365914 583018 365946 583254
rect 366182 583018 366266 583254
rect 366502 583018 366534 583254
rect 365914 547574 366534 583018
rect 365914 547338 365946 547574
rect 366182 547338 366266 547574
rect 366502 547338 366534 547574
rect 365914 547254 366534 547338
rect 365914 547018 365946 547254
rect 366182 547018 366266 547254
rect 366502 547018 366534 547254
rect 365914 511574 366534 547018
rect 365914 511338 365946 511574
rect 366182 511338 366266 511574
rect 366502 511338 366534 511574
rect 365914 511254 366534 511338
rect 365914 511018 365946 511254
rect 366182 511018 366266 511254
rect 366502 511018 366534 511254
rect 365914 475574 366534 511018
rect 365914 475338 365946 475574
rect 366182 475338 366266 475574
rect 366502 475338 366534 475574
rect 365914 475254 366534 475338
rect 365914 475018 365946 475254
rect 366182 475018 366266 475254
rect 366502 475018 366534 475254
rect 365914 439574 366534 475018
rect 365914 439338 365946 439574
rect 366182 439338 366266 439574
rect 366502 439338 366534 439574
rect 365914 439254 366534 439338
rect 365914 439018 365946 439254
rect 366182 439018 366266 439254
rect 366502 439018 366534 439254
rect 365914 403574 366534 439018
rect 365914 403338 365946 403574
rect 366182 403338 366266 403574
rect 366502 403338 366534 403574
rect 365914 403254 366534 403338
rect 365914 403018 365946 403254
rect 366182 403018 366266 403254
rect 366502 403018 366534 403254
rect 365914 367574 366534 403018
rect 365914 367338 365946 367574
rect 366182 367338 366266 367574
rect 366502 367338 366534 367574
rect 365914 367254 366534 367338
rect 365914 367018 365946 367254
rect 366182 367018 366266 367254
rect 366502 367018 366534 367254
rect 365914 331574 366534 367018
rect 365914 331338 365946 331574
rect 366182 331338 366266 331574
rect 366502 331338 366534 331574
rect 365914 331254 366534 331338
rect 365914 331018 365946 331254
rect 366182 331018 366266 331254
rect 366502 331018 366534 331254
rect 365914 295574 366534 331018
rect 365914 295338 365946 295574
rect 366182 295338 366266 295574
rect 366502 295338 366534 295574
rect 365914 295254 366534 295338
rect 365914 295018 365946 295254
rect 366182 295018 366266 295254
rect 366502 295018 366534 295254
rect 365914 259574 366534 295018
rect 365914 259338 365946 259574
rect 366182 259338 366266 259574
rect 366502 259338 366534 259574
rect 365914 259254 366534 259338
rect 365914 259018 365946 259254
rect 366182 259018 366266 259254
rect 366502 259018 366534 259254
rect 365914 223574 366534 259018
rect 365914 223338 365946 223574
rect 366182 223338 366266 223574
rect 366502 223338 366534 223574
rect 365914 223254 366534 223338
rect 365914 223018 365946 223254
rect 366182 223018 366266 223254
rect 366502 223018 366534 223254
rect 365914 187574 366534 223018
rect 365914 187338 365946 187574
rect 366182 187338 366266 187574
rect 366502 187338 366534 187574
rect 365914 187254 366534 187338
rect 365914 187018 365946 187254
rect 366182 187018 366266 187254
rect 366502 187018 366534 187254
rect 365914 151574 366534 187018
rect 365914 151338 365946 151574
rect 366182 151338 366266 151574
rect 366502 151338 366534 151574
rect 365914 151254 366534 151338
rect 365914 151018 365946 151254
rect 366182 151018 366266 151254
rect 366502 151018 366534 151254
rect 365914 115574 366534 151018
rect 365914 115338 365946 115574
rect 366182 115338 366266 115574
rect 366502 115338 366534 115574
rect 365914 115254 366534 115338
rect 365914 115018 365946 115254
rect 366182 115018 366266 115254
rect 366502 115018 366534 115254
rect 365914 79574 366534 115018
rect 365914 79338 365946 79574
rect 366182 79338 366266 79574
rect 366502 79338 366534 79574
rect 365914 79254 366534 79338
rect 365914 79018 365946 79254
rect 366182 79018 366266 79254
rect 366502 79018 366534 79254
rect 365914 43574 366534 79018
rect 365914 43338 365946 43574
rect 366182 43338 366266 43574
rect 366502 43338 366534 43574
rect 365914 43254 366534 43338
rect 365914 43018 365946 43254
rect 366182 43018 366266 43254
rect 366502 43018 366534 43254
rect 365914 7574 366534 43018
rect 365914 7338 365946 7574
rect 366182 7338 366266 7574
rect 366502 7338 366534 7574
rect 365914 7254 366534 7338
rect 365914 7018 365946 7254
rect 366182 7018 366266 7254
rect 366502 7018 366534 7254
rect 365914 -1306 366534 7018
rect 365914 -1542 365946 -1306
rect 366182 -1542 366266 -1306
rect 366502 -1542 366534 -1306
rect 365914 -1626 366534 -1542
rect 365914 -1862 365946 -1626
rect 366182 -1862 366266 -1626
rect 366502 -1862 366534 -1626
rect 365914 -7654 366534 -1862
rect 369634 706758 370254 711590
rect 369634 706522 369666 706758
rect 369902 706522 369986 706758
rect 370222 706522 370254 706758
rect 369634 706438 370254 706522
rect 369634 706202 369666 706438
rect 369902 706202 369986 706438
rect 370222 706202 370254 706438
rect 369634 695294 370254 706202
rect 369634 695058 369666 695294
rect 369902 695058 369986 695294
rect 370222 695058 370254 695294
rect 369634 694974 370254 695058
rect 369634 694738 369666 694974
rect 369902 694738 369986 694974
rect 370222 694738 370254 694974
rect 369634 659294 370254 694738
rect 369634 659058 369666 659294
rect 369902 659058 369986 659294
rect 370222 659058 370254 659294
rect 369634 658974 370254 659058
rect 369634 658738 369666 658974
rect 369902 658738 369986 658974
rect 370222 658738 370254 658974
rect 369634 623294 370254 658738
rect 369634 623058 369666 623294
rect 369902 623058 369986 623294
rect 370222 623058 370254 623294
rect 369634 622974 370254 623058
rect 369634 622738 369666 622974
rect 369902 622738 369986 622974
rect 370222 622738 370254 622974
rect 369634 587294 370254 622738
rect 369634 587058 369666 587294
rect 369902 587058 369986 587294
rect 370222 587058 370254 587294
rect 369634 586974 370254 587058
rect 369634 586738 369666 586974
rect 369902 586738 369986 586974
rect 370222 586738 370254 586974
rect 369634 551294 370254 586738
rect 369634 551058 369666 551294
rect 369902 551058 369986 551294
rect 370222 551058 370254 551294
rect 369634 550974 370254 551058
rect 369634 550738 369666 550974
rect 369902 550738 369986 550974
rect 370222 550738 370254 550974
rect 369634 515294 370254 550738
rect 369634 515058 369666 515294
rect 369902 515058 369986 515294
rect 370222 515058 370254 515294
rect 369634 514974 370254 515058
rect 369634 514738 369666 514974
rect 369902 514738 369986 514974
rect 370222 514738 370254 514974
rect 369634 479294 370254 514738
rect 369634 479058 369666 479294
rect 369902 479058 369986 479294
rect 370222 479058 370254 479294
rect 369634 478974 370254 479058
rect 369634 478738 369666 478974
rect 369902 478738 369986 478974
rect 370222 478738 370254 478974
rect 369634 443294 370254 478738
rect 369634 443058 369666 443294
rect 369902 443058 369986 443294
rect 370222 443058 370254 443294
rect 369634 442974 370254 443058
rect 369634 442738 369666 442974
rect 369902 442738 369986 442974
rect 370222 442738 370254 442974
rect 369634 407294 370254 442738
rect 369634 407058 369666 407294
rect 369902 407058 369986 407294
rect 370222 407058 370254 407294
rect 369634 406974 370254 407058
rect 369634 406738 369666 406974
rect 369902 406738 369986 406974
rect 370222 406738 370254 406974
rect 369634 371294 370254 406738
rect 369634 371058 369666 371294
rect 369902 371058 369986 371294
rect 370222 371058 370254 371294
rect 369634 370974 370254 371058
rect 369634 370738 369666 370974
rect 369902 370738 369986 370974
rect 370222 370738 370254 370974
rect 369634 335294 370254 370738
rect 369634 335058 369666 335294
rect 369902 335058 369986 335294
rect 370222 335058 370254 335294
rect 369634 334974 370254 335058
rect 369634 334738 369666 334974
rect 369902 334738 369986 334974
rect 370222 334738 370254 334974
rect 369634 299294 370254 334738
rect 369634 299058 369666 299294
rect 369902 299058 369986 299294
rect 370222 299058 370254 299294
rect 369634 298974 370254 299058
rect 369634 298738 369666 298974
rect 369902 298738 369986 298974
rect 370222 298738 370254 298974
rect 369634 263294 370254 298738
rect 369634 263058 369666 263294
rect 369902 263058 369986 263294
rect 370222 263058 370254 263294
rect 369634 262974 370254 263058
rect 369634 262738 369666 262974
rect 369902 262738 369986 262974
rect 370222 262738 370254 262974
rect 369634 227294 370254 262738
rect 369634 227058 369666 227294
rect 369902 227058 369986 227294
rect 370222 227058 370254 227294
rect 369634 226974 370254 227058
rect 369634 226738 369666 226974
rect 369902 226738 369986 226974
rect 370222 226738 370254 226974
rect 369634 191294 370254 226738
rect 369634 191058 369666 191294
rect 369902 191058 369986 191294
rect 370222 191058 370254 191294
rect 369634 190974 370254 191058
rect 369634 190738 369666 190974
rect 369902 190738 369986 190974
rect 370222 190738 370254 190974
rect 369634 155294 370254 190738
rect 369634 155058 369666 155294
rect 369902 155058 369986 155294
rect 370222 155058 370254 155294
rect 369634 154974 370254 155058
rect 369634 154738 369666 154974
rect 369902 154738 369986 154974
rect 370222 154738 370254 154974
rect 369634 119294 370254 154738
rect 369634 119058 369666 119294
rect 369902 119058 369986 119294
rect 370222 119058 370254 119294
rect 369634 118974 370254 119058
rect 369634 118738 369666 118974
rect 369902 118738 369986 118974
rect 370222 118738 370254 118974
rect 369634 83294 370254 118738
rect 369634 83058 369666 83294
rect 369902 83058 369986 83294
rect 370222 83058 370254 83294
rect 369634 82974 370254 83058
rect 369634 82738 369666 82974
rect 369902 82738 369986 82974
rect 370222 82738 370254 82974
rect 369634 47294 370254 82738
rect 369634 47058 369666 47294
rect 369902 47058 369986 47294
rect 370222 47058 370254 47294
rect 369634 46974 370254 47058
rect 369634 46738 369666 46974
rect 369902 46738 369986 46974
rect 370222 46738 370254 46974
rect 369634 11294 370254 46738
rect 369634 11058 369666 11294
rect 369902 11058 369986 11294
rect 370222 11058 370254 11294
rect 369634 10974 370254 11058
rect 369634 10738 369666 10974
rect 369902 10738 369986 10974
rect 370222 10738 370254 10974
rect 369634 -2266 370254 10738
rect 369634 -2502 369666 -2266
rect 369902 -2502 369986 -2266
rect 370222 -2502 370254 -2266
rect 369634 -2586 370254 -2502
rect 369634 -2822 369666 -2586
rect 369902 -2822 369986 -2586
rect 370222 -2822 370254 -2586
rect 369634 -7654 370254 -2822
rect 373354 707718 373974 711590
rect 373354 707482 373386 707718
rect 373622 707482 373706 707718
rect 373942 707482 373974 707718
rect 373354 707398 373974 707482
rect 373354 707162 373386 707398
rect 373622 707162 373706 707398
rect 373942 707162 373974 707398
rect 373354 699014 373974 707162
rect 373354 698778 373386 699014
rect 373622 698778 373706 699014
rect 373942 698778 373974 699014
rect 373354 698694 373974 698778
rect 373354 698458 373386 698694
rect 373622 698458 373706 698694
rect 373942 698458 373974 698694
rect 373354 663014 373974 698458
rect 373354 662778 373386 663014
rect 373622 662778 373706 663014
rect 373942 662778 373974 663014
rect 373354 662694 373974 662778
rect 373354 662458 373386 662694
rect 373622 662458 373706 662694
rect 373942 662458 373974 662694
rect 373354 627014 373974 662458
rect 373354 626778 373386 627014
rect 373622 626778 373706 627014
rect 373942 626778 373974 627014
rect 373354 626694 373974 626778
rect 373354 626458 373386 626694
rect 373622 626458 373706 626694
rect 373942 626458 373974 626694
rect 373354 591014 373974 626458
rect 373354 590778 373386 591014
rect 373622 590778 373706 591014
rect 373942 590778 373974 591014
rect 373354 590694 373974 590778
rect 373354 590458 373386 590694
rect 373622 590458 373706 590694
rect 373942 590458 373974 590694
rect 373354 555014 373974 590458
rect 373354 554778 373386 555014
rect 373622 554778 373706 555014
rect 373942 554778 373974 555014
rect 373354 554694 373974 554778
rect 373354 554458 373386 554694
rect 373622 554458 373706 554694
rect 373942 554458 373974 554694
rect 373354 519014 373974 554458
rect 373354 518778 373386 519014
rect 373622 518778 373706 519014
rect 373942 518778 373974 519014
rect 373354 518694 373974 518778
rect 373354 518458 373386 518694
rect 373622 518458 373706 518694
rect 373942 518458 373974 518694
rect 373354 483014 373974 518458
rect 373354 482778 373386 483014
rect 373622 482778 373706 483014
rect 373942 482778 373974 483014
rect 373354 482694 373974 482778
rect 373354 482458 373386 482694
rect 373622 482458 373706 482694
rect 373942 482458 373974 482694
rect 373354 447014 373974 482458
rect 373354 446778 373386 447014
rect 373622 446778 373706 447014
rect 373942 446778 373974 447014
rect 373354 446694 373974 446778
rect 373354 446458 373386 446694
rect 373622 446458 373706 446694
rect 373942 446458 373974 446694
rect 373354 411014 373974 446458
rect 373354 410778 373386 411014
rect 373622 410778 373706 411014
rect 373942 410778 373974 411014
rect 373354 410694 373974 410778
rect 373354 410458 373386 410694
rect 373622 410458 373706 410694
rect 373942 410458 373974 410694
rect 373354 375014 373974 410458
rect 373354 374778 373386 375014
rect 373622 374778 373706 375014
rect 373942 374778 373974 375014
rect 373354 374694 373974 374778
rect 373354 374458 373386 374694
rect 373622 374458 373706 374694
rect 373942 374458 373974 374694
rect 373354 339014 373974 374458
rect 373354 338778 373386 339014
rect 373622 338778 373706 339014
rect 373942 338778 373974 339014
rect 373354 338694 373974 338778
rect 373354 338458 373386 338694
rect 373622 338458 373706 338694
rect 373942 338458 373974 338694
rect 373354 303014 373974 338458
rect 373354 302778 373386 303014
rect 373622 302778 373706 303014
rect 373942 302778 373974 303014
rect 373354 302694 373974 302778
rect 373354 302458 373386 302694
rect 373622 302458 373706 302694
rect 373942 302458 373974 302694
rect 373354 267014 373974 302458
rect 373354 266778 373386 267014
rect 373622 266778 373706 267014
rect 373942 266778 373974 267014
rect 373354 266694 373974 266778
rect 373354 266458 373386 266694
rect 373622 266458 373706 266694
rect 373942 266458 373974 266694
rect 373354 231014 373974 266458
rect 373354 230778 373386 231014
rect 373622 230778 373706 231014
rect 373942 230778 373974 231014
rect 373354 230694 373974 230778
rect 373354 230458 373386 230694
rect 373622 230458 373706 230694
rect 373942 230458 373974 230694
rect 373354 195014 373974 230458
rect 373354 194778 373386 195014
rect 373622 194778 373706 195014
rect 373942 194778 373974 195014
rect 373354 194694 373974 194778
rect 373354 194458 373386 194694
rect 373622 194458 373706 194694
rect 373942 194458 373974 194694
rect 373354 159014 373974 194458
rect 373354 158778 373386 159014
rect 373622 158778 373706 159014
rect 373942 158778 373974 159014
rect 373354 158694 373974 158778
rect 373354 158458 373386 158694
rect 373622 158458 373706 158694
rect 373942 158458 373974 158694
rect 373354 123014 373974 158458
rect 373354 122778 373386 123014
rect 373622 122778 373706 123014
rect 373942 122778 373974 123014
rect 373354 122694 373974 122778
rect 373354 122458 373386 122694
rect 373622 122458 373706 122694
rect 373942 122458 373974 122694
rect 373354 87014 373974 122458
rect 373354 86778 373386 87014
rect 373622 86778 373706 87014
rect 373942 86778 373974 87014
rect 373354 86694 373974 86778
rect 373354 86458 373386 86694
rect 373622 86458 373706 86694
rect 373942 86458 373974 86694
rect 373354 51014 373974 86458
rect 373354 50778 373386 51014
rect 373622 50778 373706 51014
rect 373942 50778 373974 51014
rect 373354 50694 373974 50778
rect 373354 50458 373386 50694
rect 373622 50458 373706 50694
rect 373942 50458 373974 50694
rect 373354 15014 373974 50458
rect 373354 14778 373386 15014
rect 373622 14778 373706 15014
rect 373942 14778 373974 15014
rect 373354 14694 373974 14778
rect 373354 14458 373386 14694
rect 373622 14458 373706 14694
rect 373942 14458 373974 14694
rect 373354 -3226 373974 14458
rect 373354 -3462 373386 -3226
rect 373622 -3462 373706 -3226
rect 373942 -3462 373974 -3226
rect 373354 -3546 373974 -3462
rect 373354 -3782 373386 -3546
rect 373622 -3782 373706 -3546
rect 373942 -3782 373974 -3546
rect 373354 -7654 373974 -3782
rect 377074 708678 377694 711590
rect 377074 708442 377106 708678
rect 377342 708442 377426 708678
rect 377662 708442 377694 708678
rect 377074 708358 377694 708442
rect 377074 708122 377106 708358
rect 377342 708122 377426 708358
rect 377662 708122 377694 708358
rect 377074 666734 377694 708122
rect 377074 666498 377106 666734
rect 377342 666498 377426 666734
rect 377662 666498 377694 666734
rect 377074 666414 377694 666498
rect 377074 666178 377106 666414
rect 377342 666178 377426 666414
rect 377662 666178 377694 666414
rect 377074 630734 377694 666178
rect 377074 630498 377106 630734
rect 377342 630498 377426 630734
rect 377662 630498 377694 630734
rect 377074 630414 377694 630498
rect 377074 630178 377106 630414
rect 377342 630178 377426 630414
rect 377662 630178 377694 630414
rect 377074 594734 377694 630178
rect 377074 594498 377106 594734
rect 377342 594498 377426 594734
rect 377662 594498 377694 594734
rect 377074 594414 377694 594498
rect 377074 594178 377106 594414
rect 377342 594178 377426 594414
rect 377662 594178 377694 594414
rect 377074 558734 377694 594178
rect 377074 558498 377106 558734
rect 377342 558498 377426 558734
rect 377662 558498 377694 558734
rect 377074 558414 377694 558498
rect 377074 558178 377106 558414
rect 377342 558178 377426 558414
rect 377662 558178 377694 558414
rect 377074 522734 377694 558178
rect 377074 522498 377106 522734
rect 377342 522498 377426 522734
rect 377662 522498 377694 522734
rect 377074 522414 377694 522498
rect 377074 522178 377106 522414
rect 377342 522178 377426 522414
rect 377662 522178 377694 522414
rect 377074 486734 377694 522178
rect 377074 486498 377106 486734
rect 377342 486498 377426 486734
rect 377662 486498 377694 486734
rect 377074 486414 377694 486498
rect 377074 486178 377106 486414
rect 377342 486178 377426 486414
rect 377662 486178 377694 486414
rect 377074 450734 377694 486178
rect 377074 450498 377106 450734
rect 377342 450498 377426 450734
rect 377662 450498 377694 450734
rect 377074 450414 377694 450498
rect 377074 450178 377106 450414
rect 377342 450178 377426 450414
rect 377662 450178 377694 450414
rect 377074 414734 377694 450178
rect 377074 414498 377106 414734
rect 377342 414498 377426 414734
rect 377662 414498 377694 414734
rect 377074 414414 377694 414498
rect 377074 414178 377106 414414
rect 377342 414178 377426 414414
rect 377662 414178 377694 414414
rect 377074 378734 377694 414178
rect 377074 378498 377106 378734
rect 377342 378498 377426 378734
rect 377662 378498 377694 378734
rect 377074 378414 377694 378498
rect 377074 378178 377106 378414
rect 377342 378178 377426 378414
rect 377662 378178 377694 378414
rect 377074 342734 377694 378178
rect 377074 342498 377106 342734
rect 377342 342498 377426 342734
rect 377662 342498 377694 342734
rect 377074 342414 377694 342498
rect 377074 342178 377106 342414
rect 377342 342178 377426 342414
rect 377662 342178 377694 342414
rect 377074 306734 377694 342178
rect 377074 306498 377106 306734
rect 377342 306498 377426 306734
rect 377662 306498 377694 306734
rect 377074 306414 377694 306498
rect 377074 306178 377106 306414
rect 377342 306178 377426 306414
rect 377662 306178 377694 306414
rect 377074 270734 377694 306178
rect 377074 270498 377106 270734
rect 377342 270498 377426 270734
rect 377662 270498 377694 270734
rect 377074 270414 377694 270498
rect 377074 270178 377106 270414
rect 377342 270178 377426 270414
rect 377662 270178 377694 270414
rect 377074 234734 377694 270178
rect 377074 234498 377106 234734
rect 377342 234498 377426 234734
rect 377662 234498 377694 234734
rect 377074 234414 377694 234498
rect 377074 234178 377106 234414
rect 377342 234178 377426 234414
rect 377662 234178 377694 234414
rect 377074 198734 377694 234178
rect 377074 198498 377106 198734
rect 377342 198498 377426 198734
rect 377662 198498 377694 198734
rect 377074 198414 377694 198498
rect 377074 198178 377106 198414
rect 377342 198178 377426 198414
rect 377662 198178 377694 198414
rect 377074 162734 377694 198178
rect 377074 162498 377106 162734
rect 377342 162498 377426 162734
rect 377662 162498 377694 162734
rect 377074 162414 377694 162498
rect 377074 162178 377106 162414
rect 377342 162178 377426 162414
rect 377662 162178 377694 162414
rect 377074 126734 377694 162178
rect 377074 126498 377106 126734
rect 377342 126498 377426 126734
rect 377662 126498 377694 126734
rect 377074 126414 377694 126498
rect 377074 126178 377106 126414
rect 377342 126178 377426 126414
rect 377662 126178 377694 126414
rect 377074 90734 377694 126178
rect 377074 90498 377106 90734
rect 377342 90498 377426 90734
rect 377662 90498 377694 90734
rect 377074 90414 377694 90498
rect 377074 90178 377106 90414
rect 377342 90178 377426 90414
rect 377662 90178 377694 90414
rect 377074 54734 377694 90178
rect 377074 54498 377106 54734
rect 377342 54498 377426 54734
rect 377662 54498 377694 54734
rect 377074 54414 377694 54498
rect 377074 54178 377106 54414
rect 377342 54178 377426 54414
rect 377662 54178 377694 54414
rect 377074 18734 377694 54178
rect 377074 18498 377106 18734
rect 377342 18498 377426 18734
rect 377662 18498 377694 18734
rect 377074 18414 377694 18498
rect 377074 18178 377106 18414
rect 377342 18178 377426 18414
rect 377662 18178 377694 18414
rect 377074 -4186 377694 18178
rect 377074 -4422 377106 -4186
rect 377342 -4422 377426 -4186
rect 377662 -4422 377694 -4186
rect 377074 -4506 377694 -4422
rect 377074 -4742 377106 -4506
rect 377342 -4742 377426 -4506
rect 377662 -4742 377694 -4506
rect 377074 -7654 377694 -4742
rect 380794 709638 381414 711590
rect 380794 709402 380826 709638
rect 381062 709402 381146 709638
rect 381382 709402 381414 709638
rect 380794 709318 381414 709402
rect 380794 709082 380826 709318
rect 381062 709082 381146 709318
rect 381382 709082 381414 709318
rect 380794 670454 381414 709082
rect 380794 670218 380826 670454
rect 381062 670218 381146 670454
rect 381382 670218 381414 670454
rect 380794 670134 381414 670218
rect 380794 669898 380826 670134
rect 381062 669898 381146 670134
rect 381382 669898 381414 670134
rect 380794 634454 381414 669898
rect 380794 634218 380826 634454
rect 381062 634218 381146 634454
rect 381382 634218 381414 634454
rect 380794 634134 381414 634218
rect 380794 633898 380826 634134
rect 381062 633898 381146 634134
rect 381382 633898 381414 634134
rect 380794 598454 381414 633898
rect 380794 598218 380826 598454
rect 381062 598218 381146 598454
rect 381382 598218 381414 598454
rect 380794 598134 381414 598218
rect 380794 597898 380826 598134
rect 381062 597898 381146 598134
rect 381382 597898 381414 598134
rect 380794 562454 381414 597898
rect 380794 562218 380826 562454
rect 381062 562218 381146 562454
rect 381382 562218 381414 562454
rect 380794 562134 381414 562218
rect 380794 561898 380826 562134
rect 381062 561898 381146 562134
rect 381382 561898 381414 562134
rect 380794 526454 381414 561898
rect 380794 526218 380826 526454
rect 381062 526218 381146 526454
rect 381382 526218 381414 526454
rect 380794 526134 381414 526218
rect 380794 525898 380826 526134
rect 381062 525898 381146 526134
rect 381382 525898 381414 526134
rect 380794 490454 381414 525898
rect 380794 490218 380826 490454
rect 381062 490218 381146 490454
rect 381382 490218 381414 490454
rect 380794 490134 381414 490218
rect 380794 489898 380826 490134
rect 381062 489898 381146 490134
rect 381382 489898 381414 490134
rect 380794 454454 381414 489898
rect 380794 454218 380826 454454
rect 381062 454218 381146 454454
rect 381382 454218 381414 454454
rect 380794 454134 381414 454218
rect 380794 453898 380826 454134
rect 381062 453898 381146 454134
rect 381382 453898 381414 454134
rect 380794 418454 381414 453898
rect 380794 418218 380826 418454
rect 381062 418218 381146 418454
rect 381382 418218 381414 418454
rect 380794 418134 381414 418218
rect 380794 417898 380826 418134
rect 381062 417898 381146 418134
rect 381382 417898 381414 418134
rect 380794 382454 381414 417898
rect 380794 382218 380826 382454
rect 381062 382218 381146 382454
rect 381382 382218 381414 382454
rect 380794 382134 381414 382218
rect 380794 381898 380826 382134
rect 381062 381898 381146 382134
rect 381382 381898 381414 382134
rect 380794 346454 381414 381898
rect 380794 346218 380826 346454
rect 381062 346218 381146 346454
rect 381382 346218 381414 346454
rect 380794 346134 381414 346218
rect 380794 345898 380826 346134
rect 381062 345898 381146 346134
rect 381382 345898 381414 346134
rect 380794 310454 381414 345898
rect 380794 310218 380826 310454
rect 381062 310218 381146 310454
rect 381382 310218 381414 310454
rect 380794 310134 381414 310218
rect 380794 309898 380826 310134
rect 381062 309898 381146 310134
rect 381382 309898 381414 310134
rect 380794 274454 381414 309898
rect 380794 274218 380826 274454
rect 381062 274218 381146 274454
rect 381382 274218 381414 274454
rect 380794 274134 381414 274218
rect 380794 273898 380826 274134
rect 381062 273898 381146 274134
rect 381382 273898 381414 274134
rect 380794 238454 381414 273898
rect 380794 238218 380826 238454
rect 381062 238218 381146 238454
rect 381382 238218 381414 238454
rect 380794 238134 381414 238218
rect 380794 237898 380826 238134
rect 381062 237898 381146 238134
rect 381382 237898 381414 238134
rect 380794 202454 381414 237898
rect 380794 202218 380826 202454
rect 381062 202218 381146 202454
rect 381382 202218 381414 202454
rect 380794 202134 381414 202218
rect 380794 201898 380826 202134
rect 381062 201898 381146 202134
rect 381382 201898 381414 202134
rect 380794 166454 381414 201898
rect 380794 166218 380826 166454
rect 381062 166218 381146 166454
rect 381382 166218 381414 166454
rect 380794 166134 381414 166218
rect 380794 165898 380826 166134
rect 381062 165898 381146 166134
rect 381382 165898 381414 166134
rect 380794 130454 381414 165898
rect 380794 130218 380826 130454
rect 381062 130218 381146 130454
rect 381382 130218 381414 130454
rect 380794 130134 381414 130218
rect 380794 129898 380826 130134
rect 381062 129898 381146 130134
rect 381382 129898 381414 130134
rect 380794 94454 381414 129898
rect 380794 94218 380826 94454
rect 381062 94218 381146 94454
rect 381382 94218 381414 94454
rect 380794 94134 381414 94218
rect 380794 93898 380826 94134
rect 381062 93898 381146 94134
rect 381382 93898 381414 94134
rect 380794 58454 381414 93898
rect 380794 58218 380826 58454
rect 381062 58218 381146 58454
rect 381382 58218 381414 58454
rect 380794 58134 381414 58218
rect 380794 57898 380826 58134
rect 381062 57898 381146 58134
rect 381382 57898 381414 58134
rect 380794 22454 381414 57898
rect 380794 22218 380826 22454
rect 381062 22218 381146 22454
rect 381382 22218 381414 22454
rect 380794 22134 381414 22218
rect 380794 21898 380826 22134
rect 381062 21898 381146 22134
rect 381382 21898 381414 22134
rect 380794 -5146 381414 21898
rect 380794 -5382 380826 -5146
rect 381062 -5382 381146 -5146
rect 381382 -5382 381414 -5146
rect 380794 -5466 381414 -5382
rect 380794 -5702 380826 -5466
rect 381062 -5702 381146 -5466
rect 381382 -5702 381414 -5466
rect 380794 -7654 381414 -5702
rect 384514 710598 385134 711590
rect 384514 710362 384546 710598
rect 384782 710362 384866 710598
rect 385102 710362 385134 710598
rect 384514 710278 385134 710362
rect 384514 710042 384546 710278
rect 384782 710042 384866 710278
rect 385102 710042 385134 710278
rect 384514 674174 385134 710042
rect 384514 673938 384546 674174
rect 384782 673938 384866 674174
rect 385102 673938 385134 674174
rect 384514 673854 385134 673938
rect 384514 673618 384546 673854
rect 384782 673618 384866 673854
rect 385102 673618 385134 673854
rect 384514 638174 385134 673618
rect 384514 637938 384546 638174
rect 384782 637938 384866 638174
rect 385102 637938 385134 638174
rect 384514 637854 385134 637938
rect 384514 637618 384546 637854
rect 384782 637618 384866 637854
rect 385102 637618 385134 637854
rect 384514 602174 385134 637618
rect 384514 601938 384546 602174
rect 384782 601938 384866 602174
rect 385102 601938 385134 602174
rect 384514 601854 385134 601938
rect 384514 601618 384546 601854
rect 384782 601618 384866 601854
rect 385102 601618 385134 601854
rect 384514 566174 385134 601618
rect 384514 565938 384546 566174
rect 384782 565938 384866 566174
rect 385102 565938 385134 566174
rect 384514 565854 385134 565938
rect 384514 565618 384546 565854
rect 384782 565618 384866 565854
rect 385102 565618 385134 565854
rect 384514 530174 385134 565618
rect 384514 529938 384546 530174
rect 384782 529938 384866 530174
rect 385102 529938 385134 530174
rect 384514 529854 385134 529938
rect 384514 529618 384546 529854
rect 384782 529618 384866 529854
rect 385102 529618 385134 529854
rect 384514 494174 385134 529618
rect 384514 493938 384546 494174
rect 384782 493938 384866 494174
rect 385102 493938 385134 494174
rect 384514 493854 385134 493938
rect 384514 493618 384546 493854
rect 384782 493618 384866 493854
rect 385102 493618 385134 493854
rect 384514 458174 385134 493618
rect 384514 457938 384546 458174
rect 384782 457938 384866 458174
rect 385102 457938 385134 458174
rect 384514 457854 385134 457938
rect 384514 457618 384546 457854
rect 384782 457618 384866 457854
rect 385102 457618 385134 457854
rect 384514 422174 385134 457618
rect 384514 421938 384546 422174
rect 384782 421938 384866 422174
rect 385102 421938 385134 422174
rect 384514 421854 385134 421938
rect 384514 421618 384546 421854
rect 384782 421618 384866 421854
rect 385102 421618 385134 421854
rect 384514 386174 385134 421618
rect 384514 385938 384546 386174
rect 384782 385938 384866 386174
rect 385102 385938 385134 386174
rect 384514 385854 385134 385938
rect 384514 385618 384546 385854
rect 384782 385618 384866 385854
rect 385102 385618 385134 385854
rect 384514 350174 385134 385618
rect 384514 349938 384546 350174
rect 384782 349938 384866 350174
rect 385102 349938 385134 350174
rect 384514 349854 385134 349938
rect 384514 349618 384546 349854
rect 384782 349618 384866 349854
rect 385102 349618 385134 349854
rect 384514 314174 385134 349618
rect 384514 313938 384546 314174
rect 384782 313938 384866 314174
rect 385102 313938 385134 314174
rect 384514 313854 385134 313938
rect 384514 313618 384546 313854
rect 384782 313618 384866 313854
rect 385102 313618 385134 313854
rect 384514 278174 385134 313618
rect 384514 277938 384546 278174
rect 384782 277938 384866 278174
rect 385102 277938 385134 278174
rect 384514 277854 385134 277938
rect 384514 277618 384546 277854
rect 384782 277618 384866 277854
rect 385102 277618 385134 277854
rect 384514 242174 385134 277618
rect 384514 241938 384546 242174
rect 384782 241938 384866 242174
rect 385102 241938 385134 242174
rect 384514 241854 385134 241938
rect 384514 241618 384546 241854
rect 384782 241618 384866 241854
rect 385102 241618 385134 241854
rect 384514 206174 385134 241618
rect 384514 205938 384546 206174
rect 384782 205938 384866 206174
rect 385102 205938 385134 206174
rect 384514 205854 385134 205938
rect 384514 205618 384546 205854
rect 384782 205618 384866 205854
rect 385102 205618 385134 205854
rect 384514 170174 385134 205618
rect 384514 169938 384546 170174
rect 384782 169938 384866 170174
rect 385102 169938 385134 170174
rect 384514 169854 385134 169938
rect 384514 169618 384546 169854
rect 384782 169618 384866 169854
rect 385102 169618 385134 169854
rect 384514 134174 385134 169618
rect 384514 133938 384546 134174
rect 384782 133938 384866 134174
rect 385102 133938 385134 134174
rect 384514 133854 385134 133938
rect 384514 133618 384546 133854
rect 384782 133618 384866 133854
rect 385102 133618 385134 133854
rect 384514 98174 385134 133618
rect 384514 97938 384546 98174
rect 384782 97938 384866 98174
rect 385102 97938 385134 98174
rect 384514 97854 385134 97938
rect 384514 97618 384546 97854
rect 384782 97618 384866 97854
rect 385102 97618 385134 97854
rect 384514 62174 385134 97618
rect 384514 61938 384546 62174
rect 384782 61938 384866 62174
rect 385102 61938 385134 62174
rect 384514 61854 385134 61938
rect 384514 61618 384546 61854
rect 384782 61618 384866 61854
rect 385102 61618 385134 61854
rect 384514 26174 385134 61618
rect 384514 25938 384546 26174
rect 384782 25938 384866 26174
rect 385102 25938 385134 26174
rect 384514 25854 385134 25938
rect 384514 25618 384546 25854
rect 384782 25618 384866 25854
rect 385102 25618 385134 25854
rect 384514 -6106 385134 25618
rect 384514 -6342 384546 -6106
rect 384782 -6342 384866 -6106
rect 385102 -6342 385134 -6106
rect 384514 -6426 385134 -6342
rect 384514 -6662 384546 -6426
rect 384782 -6662 384866 -6426
rect 385102 -6662 385134 -6426
rect 384514 -7654 385134 -6662
rect 388234 711558 388854 711590
rect 388234 711322 388266 711558
rect 388502 711322 388586 711558
rect 388822 711322 388854 711558
rect 388234 711238 388854 711322
rect 388234 711002 388266 711238
rect 388502 711002 388586 711238
rect 388822 711002 388854 711238
rect 388234 677894 388854 711002
rect 388234 677658 388266 677894
rect 388502 677658 388586 677894
rect 388822 677658 388854 677894
rect 388234 677574 388854 677658
rect 388234 677338 388266 677574
rect 388502 677338 388586 677574
rect 388822 677338 388854 677574
rect 388234 641894 388854 677338
rect 388234 641658 388266 641894
rect 388502 641658 388586 641894
rect 388822 641658 388854 641894
rect 388234 641574 388854 641658
rect 388234 641338 388266 641574
rect 388502 641338 388586 641574
rect 388822 641338 388854 641574
rect 388234 605894 388854 641338
rect 388234 605658 388266 605894
rect 388502 605658 388586 605894
rect 388822 605658 388854 605894
rect 388234 605574 388854 605658
rect 388234 605338 388266 605574
rect 388502 605338 388586 605574
rect 388822 605338 388854 605574
rect 388234 569894 388854 605338
rect 388234 569658 388266 569894
rect 388502 569658 388586 569894
rect 388822 569658 388854 569894
rect 388234 569574 388854 569658
rect 388234 569338 388266 569574
rect 388502 569338 388586 569574
rect 388822 569338 388854 569574
rect 388234 533894 388854 569338
rect 388234 533658 388266 533894
rect 388502 533658 388586 533894
rect 388822 533658 388854 533894
rect 388234 533574 388854 533658
rect 388234 533338 388266 533574
rect 388502 533338 388586 533574
rect 388822 533338 388854 533574
rect 388234 497894 388854 533338
rect 388234 497658 388266 497894
rect 388502 497658 388586 497894
rect 388822 497658 388854 497894
rect 388234 497574 388854 497658
rect 388234 497338 388266 497574
rect 388502 497338 388586 497574
rect 388822 497338 388854 497574
rect 388234 461894 388854 497338
rect 388234 461658 388266 461894
rect 388502 461658 388586 461894
rect 388822 461658 388854 461894
rect 388234 461574 388854 461658
rect 388234 461338 388266 461574
rect 388502 461338 388586 461574
rect 388822 461338 388854 461574
rect 388234 425894 388854 461338
rect 388234 425658 388266 425894
rect 388502 425658 388586 425894
rect 388822 425658 388854 425894
rect 388234 425574 388854 425658
rect 388234 425338 388266 425574
rect 388502 425338 388586 425574
rect 388822 425338 388854 425574
rect 388234 389894 388854 425338
rect 388234 389658 388266 389894
rect 388502 389658 388586 389894
rect 388822 389658 388854 389894
rect 388234 389574 388854 389658
rect 388234 389338 388266 389574
rect 388502 389338 388586 389574
rect 388822 389338 388854 389574
rect 388234 353894 388854 389338
rect 388234 353658 388266 353894
rect 388502 353658 388586 353894
rect 388822 353658 388854 353894
rect 388234 353574 388854 353658
rect 388234 353338 388266 353574
rect 388502 353338 388586 353574
rect 388822 353338 388854 353574
rect 388234 317894 388854 353338
rect 388234 317658 388266 317894
rect 388502 317658 388586 317894
rect 388822 317658 388854 317894
rect 388234 317574 388854 317658
rect 388234 317338 388266 317574
rect 388502 317338 388586 317574
rect 388822 317338 388854 317574
rect 388234 281894 388854 317338
rect 388234 281658 388266 281894
rect 388502 281658 388586 281894
rect 388822 281658 388854 281894
rect 388234 281574 388854 281658
rect 388234 281338 388266 281574
rect 388502 281338 388586 281574
rect 388822 281338 388854 281574
rect 388234 245894 388854 281338
rect 388234 245658 388266 245894
rect 388502 245658 388586 245894
rect 388822 245658 388854 245894
rect 388234 245574 388854 245658
rect 388234 245338 388266 245574
rect 388502 245338 388586 245574
rect 388822 245338 388854 245574
rect 388234 209894 388854 245338
rect 388234 209658 388266 209894
rect 388502 209658 388586 209894
rect 388822 209658 388854 209894
rect 388234 209574 388854 209658
rect 388234 209338 388266 209574
rect 388502 209338 388586 209574
rect 388822 209338 388854 209574
rect 388234 173894 388854 209338
rect 388234 173658 388266 173894
rect 388502 173658 388586 173894
rect 388822 173658 388854 173894
rect 388234 173574 388854 173658
rect 388234 173338 388266 173574
rect 388502 173338 388586 173574
rect 388822 173338 388854 173574
rect 388234 137894 388854 173338
rect 388234 137658 388266 137894
rect 388502 137658 388586 137894
rect 388822 137658 388854 137894
rect 388234 137574 388854 137658
rect 388234 137338 388266 137574
rect 388502 137338 388586 137574
rect 388822 137338 388854 137574
rect 388234 101894 388854 137338
rect 388234 101658 388266 101894
rect 388502 101658 388586 101894
rect 388822 101658 388854 101894
rect 388234 101574 388854 101658
rect 388234 101338 388266 101574
rect 388502 101338 388586 101574
rect 388822 101338 388854 101574
rect 388234 65894 388854 101338
rect 388234 65658 388266 65894
rect 388502 65658 388586 65894
rect 388822 65658 388854 65894
rect 388234 65574 388854 65658
rect 388234 65338 388266 65574
rect 388502 65338 388586 65574
rect 388822 65338 388854 65574
rect 388234 29894 388854 65338
rect 388234 29658 388266 29894
rect 388502 29658 388586 29894
rect 388822 29658 388854 29894
rect 388234 29574 388854 29658
rect 388234 29338 388266 29574
rect 388502 29338 388586 29574
rect 388822 29338 388854 29574
rect 388234 -7066 388854 29338
rect 388234 -7302 388266 -7066
rect 388502 -7302 388586 -7066
rect 388822 -7302 388854 -7066
rect 388234 -7386 388854 -7302
rect 388234 -7622 388266 -7386
rect 388502 -7622 388586 -7386
rect 388822 -7622 388854 -7386
rect 388234 -7654 388854 -7622
rect 398194 704838 398814 711590
rect 398194 704602 398226 704838
rect 398462 704602 398546 704838
rect 398782 704602 398814 704838
rect 398194 704518 398814 704602
rect 398194 704282 398226 704518
rect 398462 704282 398546 704518
rect 398782 704282 398814 704518
rect 398194 687854 398814 704282
rect 398194 687618 398226 687854
rect 398462 687618 398546 687854
rect 398782 687618 398814 687854
rect 398194 687534 398814 687618
rect 398194 687298 398226 687534
rect 398462 687298 398546 687534
rect 398782 687298 398814 687534
rect 398194 651854 398814 687298
rect 398194 651618 398226 651854
rect 398462 651618 398546 651854
rect 398782 651618 398814 651854
rect 398194 651534 398814 651618
rect 398194 651298 398226 651534
rect 398462 651298 398546 651534
rect 398782 651298 398814 651534
rect 398194 615854 398814 651298
rect 398194 615618 398226 615854
rect 398462 615618 398546 615854
rect 398782 615618 398814 615854
rect 398194 615534 398814 615618
rect 398194 615298 398226 615534
rect 398462 615298 398546 615534
rect 398782 615298 398814 615534
rect 398194 579854 398814 615298
rect 398194 579618 398226 579854
rect 398462 579618 398546 579854
rect 398782 579618 398814 579854
rect 398194 579534 398814 579618
rect 398194 579298 398226 579534
rect 398462 579298 398546 579534
rect 398782 579298 398814 579534
rect 398194 543854 398814 579298
rect 398194 543618 398226 543854
rect 398462 543618 398546 543854
rect 398782 543618 398814 543854
rect 398194 543534 398814 543618
rect 398194 543298 398226 543534
rect 398462 543298 398546 543534
rect 398782 543298 398814 543534
rect 398194 507854 398814 543298
rect 398194 507618 398226 507854
rect 398462 507618 398546 507854
rect 398782 507618 398814 507854
rect 398194 507534 398814 507618
rect 398194 507298 398226 507534
rect 398462 507298 398546 507534
rect 398782 507298 398814 507534
rect 398194 471854 398814 507298
rect 398194 471618 398226 471854
rect 398462 471618 398546 471854
rect 398782 471618 398814 471854
rect 398194 471534 398814 471618
rect 398194 471298 398226 471534
rect 398462 471298 398546 471534
rect 398782 471298 398814 471534
rect 398194 435854 398814 471298
rect 398194 435618 398226 435854
rect 398462 435618 398546 435854
rect 398782 435618 398814 435854
rect 398194 435534 398814 435618
rect 398194 435298 398226 435534
rect 398462 435298 398546 435534
rect 398782 435298 398814 435534
rect 398194 399854 398814 435298
rect 398194 399618 398226 399854
rect 398462 399618 398546 399854
rect 398782 399618 398814 399854
rect 398194 399534 398814 399618
rect 398194 399298 398226 399534
rect 398462 399298 398546 399534
rect 398782 399298 398814 399534
rect 398194 363854 398814 399298
rect 398194 363618 398226 363854
rect 398462 363618 398546 363854
rect 398782 363618 398814 363854
rect 398194 363534 398814 363618
rect 398194 363298 398226 363534
rect 398462 363298 398546 363534
rect 398782 363298 398814 363534
rect 398194 327854 398814 363298
rect 398194 327618 398226 327854
rect 398462 327618 398546 327854
rect 398782 327618 398814 327854
rect 398194 327534 398814 327618
rect 398194 327298 398226 327534
rect 398462 327298 398546 327534
rect 398782 327298 398814 327534
rect 398194 291854 398814 327298
rect 398194 291618 398226 291854
rect 398462 291618 398546 291854
rect 398782 291618 398814 291854
rect 398194 291534 398814 291618
rect 398194 291298 398226 291534
rect 398462 291298 398546 291534
rect 398782 291298 398814 291534
rect 398194 255854 398814 291298
rect 398194 255618 398226 255854
rect 398462 255618 398546 255854
rect 398782 255618 398814 255854
rect 398194 255534 398814 255618
rect 398194 255298 398226 255534
rect 398462 255298 398546 255534
rect 398782 255298 398814 255534
rect 398194 219854 398814 255298
rect 398194 219618 398226 219854
rect 398462 219618 398546 219854
rect 398782 219618 398814 219854
rect 398194 219534 398814 219618
rect 398194 219298 398226 219534
rect 398462 219298 398546 219534
rect 398782 219298 398814 219534
rect 398194 183854 398814 219298
rect 398194 183618 398226 183854
rect 398462 183618 398546 183854
rect 398782 183618 398814 183854
rect 398194 183534 398814 183618
rect 398194 183298 398226 183534
rect 398462 183298 398546 183534
rect 398782 183298 398814 183534
rect 398194 147854 398814 183298
rect 398194 147618 398226 147854
rect 398462 147618 398546 147854
rect 398782 147618 398814 147854
rect 398194 147534 398814 147618
rect 398194 147298 398226 147534
rect 398462 147298 398546 147534
rect 398782 147298 398814 147534
rect 398194 111854 398814 147298
rect 398194 111618 398226 111854
rect 398462 111618 398546 111854
rect 398782 111618 398814 111854
rect 398194 111534 398814 111618
rect 398194 111298 398226 111534
rect 398462 111298 398546 111534
rect 398782 111298 398814 111534
rect 398194 75854 398814 111298
rect 398194 75618 398226 75854
rect 398462 75618 398546 75854
rect 398782 75618 398814 75854
rect 398194 75534 398814 75618
rect 398194 75298 398226 75534
rect 398462 75298 398546 75534
rect 398782 75298 398814 75534
rect 398194 39854 398814 75298
rect 398194 39618 398226 39854
rect 398462 39618 398546 39854
rect 398782 39618 398814 39854
rect 398194 39534 398814 39618
rect 398194 39298 398226 39534
rect 398462 39298 398546 39534
rect 398782 39298 398814 39534
rect 398194 3854 398814 39298
rect 398194 3618 398226 3854
rect 398462 3618 398546 3854
rect 398782 3618 398814 3854
rect 398194 3534 398814 3618
rect 398194 3298 398226 3534
rect 398462 3298 398546 3534
rect 398782 3298 398814 3534
rect 398194 -346 398814 3298
rect 398194 -582 398226 -346
rect 398462 -582 398546 -346
rect 398782 -582 398814 -346
rect 398194 -666 398814 -582
rect 398194 -902 398226 -666
rect 398462 -902 398546 -666
rect 398782 -902 398814 -666
rect 398194 -7654 398814 -902
rect 401914 705798 402534 711590
rect 401914 705562 401946 705798
rect 402182 705562 402266 705798
rect 402502 705562 402534 705798
rect 401914 705478 402534 705562
rect 401914 705242 401946 705478
rect 402182 705242 402266 705478
rect 402502 705242 402534 705478
rect 401914 691574 402534 705242
rect 401914 691338 401946 691574
rect 402182 691338 402266 691574
rect 402502 691338 402534 691574
rect 401914 691254 402534 691338
rect 401914 691018 401946 691254
rect 402182 691018 402266 691254
rect 402502 691018 402534 691254
rect 401914 655574 402534 691018
rect 401914 655338 401946 655574
rect 402182 655338 402266 655574
rect 402502 655338 402534 655574
rect 401914 655254 402534 655338
rect 401914 655018 401946 655254
rect 402182 655018 402266 655254
rect 402502 655018 402534 655254
rect 401914 619574 402534 655018
rect 401914 619338 401946 619574
rect 402182 619338 402266 619574
rect 402502 619338 402534 619574
rect 401914 619254 402534 619338
rect 401914 619018 401946 619254
rect 402182 619018 402266 619254
rect 402502 619018 402534 619254
rect 401914 583574 402534 619018
rect 401914 583338 401946 583574
rect 402182 583338 402266 583574
rect 402502 583338 402534 583574
rect 401914 583254 402534 583338
rect 401914 583018 401946 583254
rect 402182 583018 402266 583254
rect 402502 583018 402534 583254
rect 401914 547574 402534 583018
rect 401914 547338 401946 547574
rect 402182 547338 402266 547574
rect 402502 547338 402534 547574
rect 401914 547254 402534 547338
rect 401914 547018 401946 547254
rect 402182 547018 402266 547254
rect 402502 547018 402534 547254
rect 401914 511574 402534 547018
rect 401914 511338 401946 511574
rect 402182 511338 402266 511574
rect 402502 511338 402534 511574
rect 401914 511254 402534 511338
rect 401914 511018 401946 511254
rect 402182 511018 402266 511254
rect 402502 511018 402534 511254
rect 401914 475574 402534 511018
rect 401914 475338 401946 475574
rect 402182 475338 402266 475574
rect 402502 475338 402534 475574
rect 401914 475254 402534 475338
rect 401914 475018 401946 475254
rect 402182 475018 402266 475254
rect 402502 475018 402534 475254
rect 401914 439574 402534 475018
rect 401914 439338 401946 439574
rect 402182 439338 402266 439574
rect 402502 439338 402534 439574
rect 401914 439254 402534 439338
rect 401914 439018 401946 439254
rect 402182 439018 402266 439254
rect 402502 439018 402534 439254
rect 401914 403574 402534 439018
rect 401914 403338 401946 403574
rect 402182 403338 402266 403574
rect 402502 403338 402534 403574
rect 401914 403254 402534 403338
rect 401914 403018 401946 403254
rect 402182 403018 402266 403254
rect 402502 403018 402534 403254
rect 401914 367574 402534 403018
rect 401914 367338 401946 367574
rect 402182 367338 402266 367574
rect 402502 367338 402534 367574
rect 401914 367254 402534 367338
rect 401914 367018 401946 367254
rect 402182 367018 402266 367254
rect 402502 367018 402534 367254
rect 401914 331574 402534 367018
rect 401914 331338 401946 331574
rect 402182 331338 402266 331574
rect 402502 331338 402534 331574
rect 401914 331254 402534 331338
rect 401914 331018 401946 331254
rect 402182 331018 402266 331254
rect 402502 331018 402534 331254
rect 401914 295574 402534 331018
rect 401914 295338 401946 295574
rect 402182 295338 402266 295574
rect 402502 295338 402534 295574
rect 401914 295254 402534 295338
rect 401914 295018 401946 295254
rect 402182 295018 402266 295254
rect 402502 295018 402534 295254
rect 401914 259574 402534 295018
rect 401914 259338 401946 259574
rect 402182 259338 402266 259574
rect 402502 259338 402534 259574
rect 401914 259254 402534 259338
rect 401914 259018 401946 259254
rect 402182 259018 402266 259254
rect 402502 259018 402534 259254
rect 401914 223574 402534 259018
rect 401914 223338 401946 223574
rect 402182 223338 402266 223574
rect 402502 223338 402534 223574
rect 401914 223254 402534 223338
rect 401914 223018 401946 223254
rect 402182 223018 402266 223254
rect 402502 223018 402534 223254
rect 401914 187574 402534 223018
rect 401914 187338 401946 187574
rect 402182 187338 402266 187574
rect 402502 187338 402534 187574
rect 401914 187254 402534 187338
rect 401914 187018 401946 187254
rect 402182 187018 402266 187254
rect 402502 187018 402534 187254
rect 401914 151574 402534 187018
rect 401914 151338 401946 151574
rect 402182 151338 402266 151574
rect 402502 151338 402534 151574
rect 401914 151254 402534 151338
rect 401914 151018 401946 151254
rect 402182 151018 402266 151254
rect 402502 151018 402534 151254
rect 401914 115574 402534 151018
rect 401914 115338 401946 115574
rect 402182 115338 402266 115574
rect 402502 115338 402534 115574
rect 401914 115254 402534 115338
rect 401914 115018 401946 115254
rect 402182 115018 402266 115254
rect 402502 115018 402534 115254
rect 401914 79574 402534 115018
rect 405634 706758 406254 711590
rect 405634 706522 405666 706758
rect 405902 706522 405986 706758
rect 406222 706522 406254 706758
rect 405634 706438 406254 706522
rect 405634 706202 405666 706438
rect 405902 706202 405986 706438
rect 406222 706202 406254 706438
rect 405634 695294 406254 706202
rect 405634 695058 405666 695294
rect 405902 695058 405986 695294
rect 406222 695058 406254 695294
rect 405634 694974 406254 695058
rect 405634 694738 405666 694974
rect 405902 694738 405986 694974
rect 406222 694738 406254 694974
rect 405634 659294 406254 694738
rect 405634 659058 405666 659294
rect 405902 659058 405986 659294
rect 406222 659058 406254 659294
rect 405634 658974 406254 659058
rect 405634 658738 405666 658974
rect 405902 658738 405986 658974
rect 406222 658738 406254 658974
rect 405634 623294 406254 658738
rect 405634 623058 405666 623294
rect 405902 623058 405986 623294
rect 406222 623058 406254 623294
rect 405634 622974 406254 623058
rect 405634 622738 405666 622974
rect 405902 622738 405986 622974
rect 406222 622738 406254 622974
rect 405634 587294 406254 622738
rect 405634 587058 405666 587294
rect 405902 587058 405986 587294
rect 406222 587058 406254 587294
rect 405634 586974 406254 587058
rect 405634 586738 405666 586974
rect 405902 586738 405986 586974
rect 406222 586738 406254 586974
rect 405634 551294 406254 586738
rect 405634 551058 405666 551294
rect 405902 551058 405986 551294
rect 406222 551058 406254 551294
rect 405634 550974 406254 551058
rect 405634 550738 405666 550974
rect 405902 550738 405986 550974
rect 406222 550738 406254 550974
rect 405634 515294 406254 550738
rect 405634 515058 405666 515294
rect 405902 515058 405986 515294
rect 406222 515058 406254 515294
rect 405634 514974 406254 515058
rect 405634 514738 405666 514974
rect 405902 514738 405986 514974
rect 406222 514738 406254 514974
rect 405634 479294 406254 514738
rect 405634 479058 405666 479294
rect 405902 479058 405986 479294
rect 406222 479058 406254 479294
rect 405634 478974 406254 479058
rect 405634 478738 405666 478974
rect 405902 478738 405986 478974
rect 406222 478738 406254 478974
rect 405634 443294 406254 478738
rect 405634 443058 405666 443294
rect 405902 443058 405986 443294
rect 406222 443058 406254 443294
rect 405634 442974 406254 443058
rect 405634 442738 405666 442974
rect 405902 442738 405986 442974
rect 406222 442738 406254 442974
rect 405634 407294 406254 442738
rect 405634 407058 405666 407294
rect 405902 407058 405986 407294
rect 406222 407058 406254 407294
rect 405634 406974 406254 407058
rect 405634 406738 405666 406974
rect 405902 406738 405986 406974
rect 406222 406738 406254 406974
rect 405634 371294 406254 406738
rect 405634 371058 405666 371294
rect 405902 371058 405986 371294
rect 406222 371058 406254 371294
rect 405634 370974 406254 371058
rect 405634 370738 405666 370974
rect 405902 370738 405986 370974
rect 406222 370738 406254 370974
rect 405634 335294 406254 370738
rect 405634 335058 405666 335294
rect 405902 335058 405986 335294
rect 406222 335058 406254 335294
rect 405634 334974 406254 335058
rect 405634 334738 405666 334974
rect 405902 334738 405986 334974
rect 406222 334738 406254 334974
rect 405634 299294 406254 334738
rect 405634 299058 405666 299294
rect 405902 299058 405986 299294
rect 406222 299058 406254 299294
rect 405634 298974 406254 299058
rect 405634 298738 405666 298974
rect 405902 298738 405986 298974
rect 406222 298738 406254 298974
rect 405634 263294 406254 298738
rect 405634 263058 405666 263294
rect 405902 263058 405986 263294
rect 406222 263058 406254 263294
rect 405634 262974 406254 263058
rect 405634 262738 405666 262974
rect 405902 262738 405986 262974
rect 406222 262738 406254 262974
rect 405634 227294 406254 262738
rect 405634 227058 405666 227294
rect 405902 227058 405986 227294
rect 406222 227058 406254 227294
rect 405634 226974 406254 227058
rect 405634 226738 405666 226974
rect 405902 226738 405986 226974
rect 406222 226738 406254 226974
rect 405634 191294 406254 226738
rect 405634 191058 405666 191294
rect 405902 191058 405986 191294
rect 406222 191058 406254 191294
rect 405634 190974 406254 191058
rect 405634 190738 405666 190974
rect 405902 190738 405986 190974
rect 406222 190738 406254 190974
rect 405634 155294 406254 190738
rect 405634 155058 405666 155294
rect 405902 155058 405986 155294
rect 406222 155058 406254 155294
rect 405634 154974 406254 155058
rect 405634 154738 405666 154974
rect 405902 154738 405986 154974
rect 406222 154738 406254 154974
rect 405634 119294 406254 154738
rect 405634 119058 405666 119294
rect 405902 119058 405986 119294
rect 406222 119058 406254 119294
rect 405634 118974 406254 119058
rect 405634 118738 405666 118974
rect 405902 118738 405986 118974
rect 406222 118738 406254 118974
rect 404208 111854 404528 111886
rect 404208 111618 404250 111854
rect 404486 111618 404528 111854
rect 404208 111534 404528 111618
rect 404208 111298 404250 111534
rect 404486 111298 404528 111534
rect 404208 111266 404528 111298
rect 401914 79338 401946 79574
rect 402182 79338 402266 79574
rect 402502 79338 402534 79574
rect 401914 79254 402534 79338
rect 401914 79018 401946 79254
rect 402182 79018 402266 79254
rect 402502 79018 402534 79254
rect 401914 43574 402534 79018
rect 401914 43338 401946 43574
rect 402182 43338 402266 43574
rect 402502 43338 402534 43574
rect 401914 43254 402534 43338
rect 401914 43018 401946 43254
rect 402182 43018 402266 43254
rect 402502 43018 402534 43254
rect 401914 7574 402534 43018
rect 401914 7338 401946 7574
rect 402182 7338 402266 7574
rect 402502 7338 402534 7574
rect 401914 7254 402534 7338
rect 401914 7018 401946 7254
rect 402182 7018 402266 7254
rect 402502 7018 402534 7254
rect 401914 -1306 402534 7018
rect 401914 -1542 401946 -1306
rect 402182 -1542 402266 -1306
rect 402502 -1542 402534 -1306
rect 401914 -1626 402534 -1542
rect 401914 -1862 401946 -1626
rect 402182 -1862 402266 -1626
rect 402502 -1862 402534 -1626
rect 401914 -7654 402534 -1862
rect 405634 83294 406254 118738
rect 405634 83058 405666 83294
rect 405902 83058 405986 83294
rect 406222 83058 406254 83294
rect 405634 82974 406254 83058
rect 405634 82738 405666 82974
rect 405902 82738 405986 82974
rect 406222 82738 406254 82974
rect 405634 47294 406254 82738
rect 409354 707718 409974 711590
rect 409354 707482 409386 707718
rect 409622 707482 409706 707718
rect 409942 707482 409974 707718
rect 409354 707398 409974 707482
rect 409354 707162 409386 707398
rect 409622 707162 409706 707398
rect 409942 707162 409974 707398
rect 409354 699014 409974 707162
rect 409354 698778 409386 699014
rect 409622 698778 409706 699014
rect 409942 698778 409974 699014
rect 409354 698694 409974 698778
rect 409354 698458 409386 698694
rect 409622 698458 409706 698694
rect 409942 698458 409974 698694
rect 409354 663014 409974 698458
rect 409354 662778 409386 663014
rect 409622 662778 409706 663014
rect 409942 662778 409974 663014
rect 409354 662694 409974 662778
rect 409354 662458 409386 662694
rect 409622 662458 409706 662694
rect 409942 662458 409974 662694
rect 409354 627014 409974 662458
rect 409354 626778 409386 627014
rect 409622 626778 409706 627014
rect 409942 626778 409974 627014
rect 409354 626694 409974 626778
rect 409354 626458 409386 626694
rect 409622 626458 409706 626694
rect 409942 626458 409974 626694
rect 409354 591014 409974 626458
rect 409354 590778 409386 591014
rect 409622 590778 409706 591014
rect 409942 590778 409974 591014
rect 409354 590694 409974 590778
rect 409354 590458 409386 590694
rect 409622 590458 409706 590694
rect 409942 590458 409974 590694
rect 409354 555014 409974 590458
rect 409354 554778 409386 555014
rect 409622 554778 409706 555014
rect 409942 554778 409974 555014
rect 409354 554694 409974 554778
rect 409354 554458 409386 554694
rect 409622 554458 409706 554694
rect 409942 554458 409974 554694
rect 409354 519014 409974 554458
rect 409354 518778 409386 519014
rect 409622 518778 409706 519014
rect 409942 518778 409974 519014
rect 409354 518694 409974 518778
rect 409354 518458 409386 518694
rect 409622 518458 409706 518694
rect 409942 518458 409974 518694
rect 409354 483014 409974 518458
rect 409354 482778 409386 483014
rect 409622 482778 409706 483014
rect 409942 482778 409974 483014
rect 409354 482694 409974 482778
rect 409354 482458 409386 482694
rect 409622 482458 409706 482694
rect 409942 482458 409974 482694
rect 409354 447014 409974 482458
rect 409354 446778 409386 447014
rect 409622 446778 409706 447014
rect 409942 446778 409974 447014
rect 409354 446694 409974 446778
rect 409354 446458 409386 446694
rect 409622 446458 409706 446694
rect 409942 446458 409974 446694
rect 409354 411014 409974 446458
rect 409354 410778 409386 411014
rect 409622 410778 409706 411014
rect 409942 410778 409974 411014
rect 409354 410694 409974 410778
rect 409354 410458 409386 410694
rect 409622 410458 409706 410694
rect 409942 410458 409974 410694
rect 409354 375014 409974 410458
rect 409354 374778 409386 375014
rect 409622 374778 409706 375014
rect 409942 374778 409974 375014
rect 409354 374694 409974 374778
rect 409354 374458 409386 374694
rect 409622 374458 409706 374694
rect 409942 374458 409974 374694
rect 409354 339014 409974 374458
rect 409354 338778 409386 339014
rect 409622 338778 409706 339014
rect 409942 338778 409974 339014
rect 409354 338694 409974 338778
rect 409354 338458 409386 338694
rect 409622 338458 409706 338694
rect 409942 338458 409974 338694
rect 409354 303014 409974 338458
rect 409354 302778 409386 303014
rect 409622 302778 409706 303014
rect 409942 302778 409974 303014
rect 409354 302694 409974 302778
rect 409354 302458 409386 302694
rect 409622 302458 409706 302694
rect 409942 302458 409974 302694
rect 409354 267014 409974 302458
rect 409354 266778 409386 267014
rect 409622 266778 409706 267014
rect 409942 266778 409974 267014
rect 409354 266694 409974 266778
rect 409354 266458 409386 266694
rect 409622 266458 409706 266694
rect 409942 266458 409974 266694
rect 409354 231014 409974 266458
rect 409354 230778 409386 231014
rect 409622 230778 409706 231014
rect 409942 230778 409974 231014
rect 409354 230694 409974 230778
rect 409354 230458 409386 230694
rect 409622 230458 409706 230694
rect 409942 230458 409974 230694
rect 409354 195014 409974 230458
rect 409354 194778 409386 195014
rect 409622 194778 409706 195014
rect 409942 194778 409974 195014
rect 409354 194694 409974 194778
rect 409354 194458 409386 194694
rect 409622 194458 409706 194694
rect 409942 194458 409974 194694
rect 409354 159014 409974 194458
rect 409354 158778 409386 159014
rect 409622 158778 409706 159014
rect 409942 158778 409974 159014
rect 409354 158694 409974 158778
rect 409354 158458 409386 158694
rect 409622 158458 409706 158694
rect 409942 158458 409974 158694
rect 409354 123014 409974 158458
rect 413074 708678 413694 711590
rect 413074 708442 413106 708678
rect 413342 708442 413426 708678
rect 413662 708442 413694 708678
rect 413074 708358 413694 708442
rect 413074 708122 413106 708358
rect 413342 708122 413426 708358
rect 413662 708122 413694 708358
rect 413074 666734 413694 708122
rect 413074 666498 413106 666734
rect 413342 666498 413426 666734
rect 413662 666498 413694 666734
rect 413074 666414 413694 666498
rect 413074 666178 413106 666414
rect 413342 666178 413426 666414
rect 413662 666178 413694 666414
rect 413074 630734 413694 666178
rect 413074 630498 413106 630734
rect 413342 630498 413426 630734
rect 413662 630498 413694 630734
rect 413074 630414 413694 630498
rect 413074 630178 413106 630414
rect 413342 630178 413426 630414
rect 413662 630178 413694 630414
rect 413074 594734 413694 630178
rect 413074 594498 413106 594734
rect 413342 594498 413426 594734
rect 413662 594498 413694 594734
rect 413074 594414 413694 594498
rect 413074 594178 413106 594414
rect 413342 594178 413426 594414
rect 413662 594178 413694 594414
rect 413074 558734 413694 594178
rect 413074 558498 413106 558734
rect 413342 558498 413426 558734
rect 413662 558498 413694 558734
rect 413074 558414 413694 558498
rect 413074 558178 413106 558414
rect 413342 558178 413426 558414
rect 413662 558178 413694 558414
rect 413074 522734 413694 558178
rect 413074 522498 413106 522734
rect 413342 522498 413426 522734
rect 413662 522498 413694 522734
rect 413074 522414 413694 522498
rect 413074 522178 413106 522414
rect 413342 522178 413426 522414
rect 413662 522178 413694 522414
rect 413074 486734 413694 522178
rect 413074 486498 413106 486734
rect 413342 486498 413426 486734
rect 413662 486498 413694 486734
rect 413074 486414 413694 486498
rect 413074 486178 413106 486414
rect 413342 486178 413426 486414
rect 413662 486178 413694 486414
rect 413074 450734 413694 486178
rect 413074 450498 413106 450734
rect 413342 450498 413426 450734
rect 413662 450498 413694 450734
rect 413074 450414 413694 450498
rect 413074 450178 413106 450414
rect 413342 450178 413426 450414
rect 413662 450178 413694 450414
rect 413074 414734 413694 450178
rect 413074 414498 413106 414734
rect 413342 414498 413426 414734
rect 413662 414498 413694 414734
rect 413074 414414 413694 414498
rect 413074 414178 413106 414414
rect 413342 414178 413426 414414
rect 413662 414178 413694 414414
rect 413074 378734 413694 414178
rect 413074 378498 413106 378734
rect 413342 378498 413426 378734
rect 413662 378498 413694 378734
rect 413074 378414 413694 378498
rect 413074 378178 413106 378414
rect 413342 378178 413426 378414
rect 413662 378178 413694 378414
rect 413074 342734 413694 378178
rect 413074 342498 413106 342734
rect 413342 342498 413426 342734
rect 413662 342498 413694 342734
rect 413074 342414 413694 342498
rect 413074 342178 413106 342414
rect 413342 342178 413426 342414
rect 413662 342178 413694 342414
rect 413074 306734 413694 342178
rect 413074 306498 413106 306734
rect 413342 306498 413426 306734
rect 413662 306498 413694 306734
rect 413074 306414 413694 306498
rect 413074 306178 413106 306414
rect 413342 306178 413426 306414
rect 413662 306178 413694 306414
rect 413074 270734 413694 306178
rect 413074 270498 413106 270734
rect 413342 270498 413426 270734
rect 413662 270498 413694 270734
rect 413074 270414 413694 270498
rect 413074 270178 413106 270414
rect 413342 270178 413426 270414
rect 413662 270178 413694 270414
rect 413074 234734 413694 270178
rect 413074 234498 413106 234734
rect 413342 234498 413426 234734
rect 413662 234498 413694 234734
rect 413074 234414 413694 234498
rect 413074 234178 413106 234414
rect 413342 234178 413426 234414
rect 413662 234178 413694 234414
rect 413074 198734 413694 234178
rect 413074 198498 413106 198734
rect 413342 198498 413426 198734
rect 413662 198498 413694 198734
rect 413074 198414 413694 198498
rect 413074 198178 413106 198414
rect 413342 198178 413426 198414
rect 413662 198178 413694 198414
rect 413074 162734 413694 198178
rect 413074 162498 413106 162734
rect 413342 162498 413426 162734
rect 413662 162498 413694 162734
rect 413074 162414 413694 162498
rect 413074 162178 413106 162414
rect 413342 162178 413426 162414
rect 413662 162178 413694 162414
rect 413074 133649 413694 162178
rect 416794 709638 417414 711590
rect 416794 709402 416826 709638
rect 417062 709402 417146 709638
rect 417382 709402 417414 709638
rect 416794 709318 417414 709402
rect 416794 709082 416826 709318
rect 417062 709082 417146 709318
rect 417382 709082 417414 709318
rect 416794 670454 417414 709082
rect 416794 670218 416826 670454
rect 417062 670218 417146 670454
rect 417382 670218 417414 670454
rect 416794 670134 417414 670218
rect 416794 669898 416826 670134
rect 417062 669898 417146 670134
rect 417382 669898 417414 670134
rect 416794 634454 417414 669898
rect 416794 634218 416826 634454
rect 417062 634218 417146 634454
rect 417382 634218 417414 634454
rect 416794 634134 417414 634218
rect 416794 633898 416826 634134
rect 417062 633898 417146 634134
rect 417382 633898 417414 634134
rect 416794 598454 417414 633898
rect 416794 598218 416826 598454
rect 417062 598218 417146 598454
rect 417382 598218 417414 598454
rect 416794 598134 417414 598218
rect 416794 597898 416826 598134
rect 417062 597898 417146 598134
rect 417382 597898 417414 598134
rect 416794 562454 417414 597898
rect 416794 562218 416826 562454
rect 417062 562218 417146 562454
rect 417382 562218 417414 562454
rect 416794 562134 417414 562218
rect 416794 561898 416826 562134
rect 417062 561898 417146 562134
rect 417382 561898 417414 562134
rect 416794 526454 417414 561898
rect 416794 526218 416826 526454
rect 417062 526218 417146 526454
rect 417382 526218 417414 526454
rect 416794 526134 417414 526218
rect 416794 525898 416826 526134
rect 417062 525898 417146 526134
rect 417382 525898 417414 526134
rect 416794 490454 417414 525898
rect 416794 490218 416826 490454
rect 417062 490218 417146 490454
rect 417382 490218 417414 490454
rect 416794 490134 417414 490218
rect 416794 489898 416826 490134
rect 417062 489898 417146 490134
rect 417382 489898 417414 490134
rect 416794 454454 417414 489898
rect 416794 454218 416826 454454
rect 417062 454218 417146 454454
rect 417382 454218 417414 454454
rect 416794 454134 417414 454218
rect 416794 453898 416826 454134
rect 417062 453898 417146 454134
rect 417382 453898 417414 454134
rect 416794 418454 417414 453898
rect 416794 418218 416826 418454
rect 417062 418218 417146 418454
rect 417382 418218 417414 418454
rect 416794 418134 417414 418218
rect 416794 417898 416826 418134
rect 417062 417898 417146 418134
rect 417382 417898 417414 418134
rect 416794 382454 417414 417898
rect 416794 382218 416826 382454
rect 417062 382218 417146 382454
rect 417382 382218 417414 382454
rect 416794 382134 417414 382218
rect 416794 381898 416826 382134
rect 417062 381898 417146 382134
rect 417382 381898 417414 382134
rect 416794 346454 417414 381898
rect 416794 346218 416826 346454
rect 417062 346218 417146 346454
rect 417382 346218 417414 346454
rect 416794 346134 417414 346218
rect 416794 345898 416826 346134
rect 417062 345898 417146 346134
rect 417382 345898 417414 346134
rect 416794 310454 417414 345898
rect 416794 310218 416826 310454
rect 417062 310218 417146 310454
rect 417382 310218 417414 310454
rect 416794 310134 417414 310218
rect 416794 309898 416826 310134
rect 417062 309898 417146 310134
rect 417382 309898 417414 310134
rect 416794 274454 417414 309898
rect 416794 274218 416826 274454
rect 417062 274218 417146 274454
rect 417382 274218 417414 274454
rect 416794 274134 417414 274218
rect 416794 273898 416826 274134
rect 417062 273898 417146 274134
rect 417382 273898 417414 274134
rect 416794 238454 417414 273898
rect 416794 238218 416826 238454
rect 417062 238218 417146 238454
rect 417382 238218 417414 238454
rect 416794 238134 417414 238218
rect 416794 237898 416826 238134
rect 417062 237898 417146 238134
rect 417382 237898 417414 238134
rect 416794 202454 417414 237898
rect 416794 202218 416826 202454
rect 417062 202218 417146 202454
rect 417382 202218 417414 202454
rect 416794 202134 417414 202218
rect 416794 201898 416826 202134
rect 417062 201898 417146 202134
rect 417382 201898 417414 202134
rect 416794 166454 417414 201898
rect 416794 166218 416826 166454
rect 417062 166218 417146 166454
rect 417382 166218 417414 166454
rect 416794 166134 417414 166218
rect 416794 165898 416826 166134
rect 417062 165898 417146 166134
rect 417382 165898 417414 166134
rect 416794 133649 417414 165898
rect 420514 710598 421134 711590
rect 420514 710362 420546 710598
rect 420782 710362 420866 710598
rect 421102 710362 421134 710598
rect 420514 710278 421134 710362
rect 420514 710042 420546 710278
rect 420782 710042 420866 710278
rect 421102 710042 421134 710278
rect 420514 674174 421134 710042
rect 420514 673938 420546 674174
rect 420782 673938 420866 674174
rect 421102 673938 421134 674174
rect 420514 673854 421134 673938
rect 420514 673618 420546 673854
rect 420782 673618 420866 673854
rect 421102 673618 421134 673854
rect 420514 638174 421134 673618
rect 420514 637938 420546 638174
rect 420782 637938 420866 638174
rect 421102 637938 421134 638174
rect 420514 637854 421134 637938
rect 420514 637618 420546 637854
rect 420782 637618 420866 637854
rect 421102 637618 421134 637854
rect 420514 602174 421134 637618
rect 420514 601938 420546 602174
rect 420782 601938 420866 602174
rect 421102 601938 421134 602174
rect 420514 601854 421134 601938
rect 420514 601618 420546 601854
rect 420782 601618 420866 601854
rect 421102 601618 421134 601854
rect 420514 566174 421134 601618
rect 420514 565938 420546 566174
rect 420782 565938 420866 566174
rect 421102 565938 421134 566174
rect 420514 565854 421134 565938
rect 420514 565618 420546 565854
rect 420782 565618 420866 565854
rect 421102 565618 421134 565854
rect 420514 530174 421134 565618
rect 420514 529938 420546 530174
rect 420782 529938 420866 530174
rect 421102 529938 421134 530174
rect 420514 529854 421134 529938
rect 420514 529618 420546 529854
rect 420782 529618 420866 529854
rect 421102 529618 421134 529854
rect 420514 494174 421134 529618
rect 420514 493938 420546 494174
rect 420782 493938 420866 494174
rect 421102 493938 421134 494174
rect 420514 493854 421134 493938
rect 420514 493618 420546 493854
rect 420782 493618 420866 493854
rect 421102 493618 421134 493854
rect 420514 458174 421134 493618
rect 420514 457938 420546 458174
rect 420782 457938 420866 458174
rect 421102 457938 421134 458174
rect 420514 457854 421134 457938
rect 420514 457618 420546 457854
rect 420782 457618 420866 457854
rect 421102 457618 421134 457854
rect 420514 422174 421134 457618
rect 420514 421938 420546 422174
rect 420782 421938 420866 422174
rect 421102 421938 421134 422174
rect 420514 421854 421134 421938
rect 420514 421618 420546 421854
rect 420782 421618 420866 421854
rect 421102 421618 421134 421854
rect 420514 386174 421134 421618
rect 420514 385938 420546 386174
rect 420782 385938 420866 386174
rect 421102 385938 421134 386174
rect 420514 385854 421134 385938
rect 420514 385618 420546 385854
rect 420782 385618 420866 385854
rect 421102 385618 421134 385854
rect 420514 350174 421134 385618
rect 420514 349938 420546 350174
rect 420782 349938 420866 350174
rect 421102 349938 421134 350174
rect 420514 349854 421134 349938
rect 420514 349618 420546 349854
rect 420782 349618 420866 349854
rect 421102 349618 421134 349854
rect 420514 314174 421134 349618
rect 420514 313938 420546 314174
rect 420782 313938 420866 314174
rect 421102 313938 421134 314174
rect 420514 313854 421134 313938
rect 420514 313618 420546 313854
rect 420782 313618 420866 313854
rect 421102 313618 421134 313854
rect 420514 278174 421134 313618
rect 420514 277938 420546 278174
rect 420782 277938 420866 278174
rect 421102 277938 421134 278174
rect 420514 277854 421134 277938
rect 420514 277618 420546 277854
rect 420782 277618 420866 277854
rect 421102 277618 421134 277854
rect 420514 242174 421134 277618
rect 420514 241938 420546 242174
rect 420782 241938 420866 242174
rect 421102 241938 421134 242174
rect 420514 241854 421134 241938
rect 420514 241618 420546 241854
rect 420782 241618 420866 241854
rect 421102 241618 421134 241854
rect 420514 206174 421134 241618
rect 420514 205938 420546 206174
rect 420782 205938 420866 206174
rect 421102 205938 421134 206174
rect 420514 205854 421134 205938
rect 420514 205618 420546 205854
rect 420782 205618 420866 205854
rect 421102 205618 421134 205854
rect 420514 170174 421134 205618
rect 420514 169938 420546 170174
rect 420782 169938 420866 170174
rect 421102 169938 421134 170174
rect 420514 169854 421134 169938
rect 420514 169618 420546 169854
rect 420782 169618 420866 169854
rect 421102 169618 421134 169854
rect 420514 134174 421134 169618
rect 420514 133938 420546 134174
rect 420782 133938 420866 134174
rect 421102 133938 421134 134174
rect 420514 133854 421134 133938
rect 420514 133618 420546 133854
rect 420782 133618 420866 133854
rect 421102 133618 421134 133854
rect 424234 711558 424854 711590
rect 424234 711322 424266 711558
rect 424502 711322 424586 711558
rect 424822 711322 424854 711558
rect 424234 711238 424854 711322
rect 424234 711002 424266 711238
rect 424502 711002 424586 711238
rect 424822 711002 424854 711238
rect 424234 677894 424854 711002
rect 424234 677658 424266 677894
rect 424502 677658 424586 677894
rect 424822 677658 424854 677894
rect 424234 677574 424854 677658
rect 424234 677338 424266 677574
rect 424502 677338 424586 677574
rect 424822 677338 424854 677574
rect 424234 641894 424854 677338
rect 424234 641658 424266 641894
rect 424502 641658 424586 641894
rect 424822 641658 424854 641894
rect 424234 641574 424854 641658
rect 424234 641338 424266 641574
rect 424502 641338 424586 641574
rect 424822 641338 424854 641574
rect 424234 605894 424854 641338
rect 424234 605658 424266 605894
rect 424502 605658 424586 605894
rect 424822 605658 424854 605894
rect 424234 605574 424854 605658
rect 424234 605338 424266 605574
rect 424502 605338 424586 605574
rect 424822 605338 424854 605574
rect 424234 569894 424854 605338
rect 424234 569658 424266 569894
rect 424502 569658 424586 569894
rect 424822 569658 424854 569894
rect 424234 569574 424854 569658
rect 424234 569338 424266 569574
rect 424502 569338 424586 569574
rect 424822 569338 424854 569574
rect 424234 533894 424854 569338
rect 424234 533658 424266 533894
rect 424502 533658 424586 533894
rect 424822 533658 424854 533894
rect 424234 533574 424854 533658
rect 424234 533338 424266 533574
rect 424502 533338 424586 533574
rect 424822 533338 424854 533574
rect 424234 497894 424854 533338
rect 424234 497658 424266 497894
rect 424502 497658 424586 497894
rect 424822 497658 424854 497894
rect 424234 497574 424854 497658
rect 424234 497338 424266 497574
rect 424502 497338 424586 497574
rect 424822 497338 424854 497574
rect 424234 461894 424854 497338
rect 424234 461658 424266 461894
rect 424502 461658 424586 461894
rect 424822 461658 424854 461894
rect 424234 461574 424854 461658
rect 424234 461338 424266 461574
rect 424502 461338 424586 461574
rect 424822 461338 424854 461574
rect 424234 425894 424854 461338
rect 424234 425658 424266 425894
rect 424502 425658 424586 425894
rect 424822 425658 424854 425894
rect 424234 425574 424854 425658
rect 424234 425338 424266 425574
rect 424502 425338 424586 425574
rect 424822 425338 424854 425574
rect 424234 389894 424854 425338
rect 424234 389658 424266 389894
rect 424502 389658 424586 389894
rect 424822 389658 424854 389894
rect 424234 389574 424854 389658
rect 424234 389338 424266 389574
rect 424502 389338 424586 389574
rect 424822 389338 424854 389574
rect 424234 353894 424854 389338
rect 424234 353658 424266 353894
rect 424502 353658 424586 353894
rect 424822 353658 424854 353894
rect 424234 353574 424854 353658
rect 424234 353338 424266 353574
rect 424502 353338 424586 353574
rect 424822 353338 424854 353574
rect 424234 317894 424854 353338
rect 424234 317658 424266 317894
rect 424502 317658 424586 317894
rect 424822 317658 424854 317894
rect 424234 317574 424854 317658
rect 424234 317338 424266 317574
rect 424502 317338 424586 317574
rect 424822 317338 424854 317574
rect 424234 281894 424854 317338
rect 424234 281658 424266 281894
rect 424502 281658 424586 281894
rect 424822 281658 424854 281894
rect 424234 281574 424854 281658
rect 424234 281338 424266 281574
rect 424502 281338 424586 281574
rect 424822 281338 424854 281574
rect 424234 245894 424854 281338
rect 424234 245658 424266 245894
rect 424502 245658 424586 245894
rect 424822 245658 424854 245894
rect 424234 245574 424854 245658
rect 424234 245338 424266 245574
rect 424502 245338 424586 245574
rect 424822 245338 424854 245574
rect 424234 209894 424854 245338
rect 424234 209658 424266 209894
rect 424502 209658 424586 209894
rect 424822 209658 424854 209894
rect 424234 209574 424854 209658
rect 424234 209338 424266 209574
rect 424502 209338 424586 209574
rect 424822 209338 424854 209574
rect 424234 173894 424854 209338
rect 424234 173658 424266 173894
rect 424502 173658 424586 173894
rect 424822 173658 424854 173894
rect 424234 173574 424854 173658
rect 424234 173338 424266 173574
rect 424502 173338 424586 173574
rect 424822 173338 424854 173574
rect 424234 137894 424854 173338
rect 424234 137658 424266 137894
rect 424502 137658 424586 137894
rect 424822 137658 424854 137894
rect 424234 137574 424854 137658
rect 424234 137338 424266 137574
rect 424502 137338 424586 137574
rect 424822 137338 424854 137574
rect 424234 133649 424854 137338
rect 434194 704838 434814 711590
rect 434194 704602 434226 704838
rect 434462 704602 434546 704838
rect 434782 704602 434814 704838
rect 434194 704518 434814 704602
rect 434194 704282 434226 704518
rect 434462 704282 434546 704518
rect 434782 704282 434814 704518
rect 434194 687854 434814 704282
rect 434194 687618 434226 687854
rect 434462 687618 434546 687854
rect 434782 687618 434814 687854
rect 434194 687534 434814 687618
rect 434194 687298 434226 687534
rect 434462 687298 434546 687534
rect 434782 687298 434814 687534
rect 434194 651854 434814 687298
rect 434194 651618 434226 651854
rect 434462 651618 434546 651854
rect 434782 651618 434814 651854
rect 434194 651534 434814 651618
rect 434194 651298 434226 651534
rect 434462 651298 434546 651534
rect 434782 651298 434814 651534
rect 434194 615854 434814 651298
rect 434194 615618 434226 615854
rect 434462 615618 434546 615854
rect 434782 615618 434814 615854
rect 434194 615534 434814 615618
rect 434194 615298 434226 615534
rect 434462 615298 434546 615534
rect 434782 615298 434814 615534
rect 434194 579854 434814 615298
rect 434194 579618 434226 579854
rect 434462 579618 434546 579854
rect 434782 579618 434814 579854
rect 434194 579534 434814 579618
rect 434194 579298 434226 579534
rect 434462 579298 434546 579534
rect 434782 579298 434814 579534
rect 434194 543854 434814 579298
rect 434194 543618 434226 543854
rect 434462 543618 434546 543854
rect 434782 543618 434814 543854
rect 434194 543534 434814 543618
rect 434194 543298 434226 543534
rect 434462 543298 434546 543534
rect 434782 543298 434814 543534
rect 434194 507854 434814 543298
rect 434194 507618 434226 507854
rect 434462 507618 434546 507854
rect 434782 507618 434814 507854
rect 434194 507534 434814 507618
rect 434194 507298 434226 507534
rect 434462 507298 434546 507534
rect 434782 507298 434814 507534
rect 434194 471854 434814 507298
rect 434194 471618 434226 471854
rect 434462 471618 434546 471854
rect 434782 471618 434814 471854
rect 434194 471534 434814 471618
rect 434194 471298 434226 471534
rect 434462 471298 434546 471534
rect 434782 471298 434814 471534
rect 434194 435854 434814 471298
rect 434194 435618 434226 435854
rect 434462 435618 434546 435854
rect 434782 435618 434814 435854
rect 434194 435534 434814 435618
rect 434194 435298 434226 435534
rect 434462 435298 434546 435534
rect 434782 435298 434814 435534
rect 434194 399854 434814 435298
rect 434194 399618 434226 399854
rect 434462 399618 434546 399854
rect 434782 399618 434814 399854
rect 434194 399534 434814 399618
rect 434194 399298 434226 399534
rect 434462 399298 434546 399534
rect 434782 399298 434814 399534
rect 434194 363854 434814 399298
rect 434194 363618 434226 363854
rect 434462 363618 434546 363854
rect 434782 363618 434814 363854
rect 434194 363534 434814 363618
rect 434194 363298 434226 363534
rect 434462 363298 434546 363534
rect 434782 363298 434814 363534
rect 434194 327854 434814 363298
rect 434194 327618 434226 327854
rect 434462 327618 434546 327854
rect 434782 327618 434814 327854
rect 434194 327534 434814 327618
rect 434194 327298 434226 327534
rect 434462 327298 434546 327534
rect 434782 327298 434814 327534
rect 434194 291854 434814 327298
rect 434194 291618 434226 291854
rect 434462 291618 434546 291854
rect 434782 291618 434814 291854
rect 434194 291534 434814 291618
rect 434194 291298 434226 291534
rect 434462 291298 434546 291534
rect 434782 291298 434814 291534
rect 434194 255854 434814 291298
rect 434194 255618 434226 255854
rect 434462 255618 434546 255854
rect 434782 255618 434814 255854
rect 434194 255534 434814 255618
rect 434194 255298 434226 255534
rect 434462 255298 434546 255534
rect 434782 255298 434814 255534
rect 434194 219854 434814 255298
rect 434194 219618 434226 219854
rect 434462 219618 434546 219854
rect 434782 219618 434814 219854
rect 434194 219534 434814 219618
rect 434194 219298 434226 219534
rect 434462 219298 434546 219534
rect 434782 219298 434814 219534
rect 434194 183854 434814 219298
rect 434194 183618 434226 183854
rect 434462 183618 434546 183854
rect 434782 183618 434814 183854
rect 434194 183534 434814 183618
rect 434194 183298 434226 183534
rect 434462 183298 434546 183534
rect 434782 183298 434814 183534
rect 434194 147854 434814 183298
rect 434194 147618 434226 147854
rect 434462 147618 434546 147854
rect 434782 147618 434814 147854
rect 434194 147534 434814 147618
rect 434194 147298 434226 147534
rect 434462 147298 434546 147534
rect 434782 147298 434814 147534
rect 434194 135500 434814 147298
rect 437914 705798 438534 711590
rect 437914 705562 437946 705798
rect 438182 705562 438266 705798
rect 438502 705562 438534 705798
rect 437914 705478 438534 705562
rect 437914 705242 437946 705478
rect 438182 705242 438266 705478
rect 438502 705242 438534 705478
rect 437914 691574 438534 705242
rect 437914 691338 437946 691574
rect 438182 691338 438266 691574
rect 438502 691338 438534 691574
rect 437914 691254 438534 691338
rect 437914 691018 437946 691254
rect 438182 691018 438266 691254
rect 438502 691018 438534 691254
rect 437914 655574 438534 691018
rect 437914 655338 437946 655574
rect 438182 655338 438266 655574
rect 438502 655338 438534 655574
rect 437914 655254 438534 655338
rect 437914 655018 437946 655254
rect 438182 655018 438266 655254
rect 438502 655018 438534 655254
rect 437914 619574 438534 655018
rect 437914 619338 437946 619574
rect 438182 619338 438266 619574
rect 438502 619338 438534 619574
rect 437914 619254 438534 619338
rect 437914 619018 437946 619254
rect 438182 619018 438266 619254
rect 438502 619018 438534 619254
rect 437914 583574 438534 619018
rect 437914 583338 437946 583574
rect 438182 583338 438266 583574
rect 438502 583338 438534 583574
rect 437914 583254 438534 583338
rect 437914 583018 437946 583254
rect 438182 583018 438266 583254
rect 438502 583018 438534 583254
rect 437914 547574 438534 583018
rect 437914 547338 437946 547574
rect 438182 547338 438266 547574
rect 438502 547338 438534 547574
rect 437914 547254 438534 547338
rect 437914 547018 437946 547254
rect 438182 547018 438266 547254
rect 438502 547018 438534 547254
rect 437914 511574 438534 547018
rect 437914 511338 437946 511574
rect 438182 511338 438266 511574
rect 438502 511338 438534 511574
rect 437914 511254 438534 511338
rect 437914 511018 437946 511254
rect 438182 511018 438266 511254
rect 438502 511018 438534 511254
rect 437914 475574 438534 511018
rect 437914 475338 437946 475574
rect 438182 475338 438266 475574
rect 438502 475338 438534 475574
rect 437914 475254 438534 475338
rect 437914 475018 437946 475254
rect 438182 475018 438266 475254
rect 438502 475018 438534 475254
rect 437914 439574 438534 475018
rect 437914 439338 437946 439574
rect 438182 439338 438266 439574
rect 438502 439338 438534 439574
rect 437914 439254 438534 439338
rect 437914 439018 437946 439254
rect 438182 439018 438266 439254
rect 438502 439018 438534 439254
rect 437914 403574 438534 439018
rect 437914 403338 437946 403574
rect 438182 403338 438266 403574
rect 438502 403338 438534 403574
rect 437914 403254 438534 403338
rect 437914 403018 437946 403254
rect 438182 403018 438266 403254
rect 438502 403018 438534 403254
rect 437914 367574 438534 403018
rect 437914 367338 437946 367574
rect 438182 367338 438266 367574
rect 438502 367338 438534 367574
rect 437914 367254 438534 367338
rect 437914 367018 437946 367254
rect 438182 367018 438266 367254
rect 438502 367018 438534 367254
rect 437914 331574 438534 367018
rect 437914 331338 437946 331574
rect 438182 331338 438266 331574
rect 438502 331338 438534 331574
rect 437914 331254 438534 331338
rect 437914 331018 437946 331254
rect 438182 331018 438266 331254
rect 438502 331018 438534 331254
rect 437914 295574 438534 331018
rect 437914 295338 437946 295574
rect 438182 295338 438266 295574
rect 438502 295338 438534 295574
rect 437914 295254 438534 295338
rect 437914 295018 437946 295254
rect 438182 295018 438266 295254
rect 438502 295018 438534 295254
rect 437914 259574 438534 295018
rect 437914 259338 437946 259574
rect 438182 259338 438266 259574
rect 438502 259338 438534 259574
rect 437914 259254 438534 259338
rect 437914 259018 437946 259254
rect 438182 259018 438266 259254
rect 438502 259018 438534 259254
rect 437914 223574 438534 259018
rect 437914 223338 437946 223574
rect 438182 223338 438266 223574
rect 438502 223338 438534 223574
rect 437914 223254 438534 223338
rect 437914 223018 437946 223254
rect 438182 223018 438266 223254
rect 438502 223018 438534 223254
rect 437914 187574 438534 223018
rect 437914 187338 437946 187574
rect 438182 187338 438266 187574
rect 438502 187338 438534 187574
rect 437914 187254 438534 187338
rect 437914 187018 437946 187254
rect 438182 187018 438266 187254
rect 438502 187018 438534 187254
rect 437914 151574 438534 187018
rect 437914 151338 437946 151574
rect 438182 151338 438266 151574
rect 438502 151338 438534 151574
rect 437914 151254 438534 151338
rect 437914 151018 437946 151254
rect 438182 151018 438266 151254
rect 438502 151018 438534 151254
rect 437914 133649 438534 151018
rect 441634 706758 442254 711590
rect 441634 706522 441666 706758
rect 441902 706522 441986 706758
rect 442222 706522 442254 706758
rect 441634 706438 442254 706522
rect 441634 706202 441666 706438
rect 441902 706202 441986 706438
rect 442222 706202 442254 706438
rect 441634 695294 442254 706202
rect 441634 695058 441666 695294
rect 441902 695058 441986 695294
rect 442222 695058 442254 695294
rect 441634 694974 442254 695058
rect 441634 694738 441666 694974
rect 441902 694738 441986 694974
rect 442222 694738 442254 694974
rect 441634 659294 442254 694738
rect 441634 659058 441666 659294
rect 441902 659058 441986 659294
rect 442222 659058 442254 659294
rect 441634 658974 442254 659058
rect 441634 658738 441666 658974
rect 441902 658738 441986 658974
rect 442222 658738 442254 658974
rect 441634 623294 442254 658738
rect 441634 623058 441666 623294
rect 441902 623058 441986 623294
rect 442222 623058 442254 623294
rect 441634 622974 442254 623058
rect 441634 622738 441666 622974
rect 441902 622738 441986 622974
rect 442222 622738 442254 622974
rect 441634 587294 442254 622738
rect 441634 587058 441666 587294
rect 441902 587058 441986 587294
rect 442222 587058 442254 587294
rect 441634 586974 442254 587058
rect 441634 586738 441666 586974
rect 441902 586738 441986 586974
rect 442222 586738 442254 586974
rect 441634 551294 442254 586738
rect 441634 551058 441666 551294
rect 441902 551058 441986 551294
rect 442222 551058 442254 551294
rect 441634 550974 442254 551058
rect 441634 550738 441666 550974
rect 441902 550738 441986 550974
rect 442222 550738 442254 550974
rect 441634 515294 442254 550738
rect 441634 515058 441666 515294
rect 441902 515058 441986 515294
rect 442222 515058 442254 515294
rect 441634 514974 442254 515058
rect 441634 514738 441666 514974
rect 441902 514738 441986 514974
rect 442222 514738 442254 514974
rect 441634 479294 442254 514738
rect 441634 479058 441666 479294
rect 441902 479058 441986 479294
rect 442222 479058 442254 479294
rect 441634 478974 442254 479058
rect 441634 478738 441666 478974
rect 441902 478738 441986 478974
rect 442222 478738 442254 478974
rect 441634 443294 442254 478738
rect 441634 443058 441666 443294
rect 441902 443058 441986 443294
rect 442222 443058 442254 443294
rect 441634 442974 442254 443058
rect 441634 442738 441666 442974
rect 441902 442738 441986 442974
rect 442222 442738 442254 442974
rect 441634 407294 442254 442738
rect 441634 407058 441666 407294
rect 441902 407058 441986 407294
rect 442222 407058 442254 407294
rect 441634 406974 442254 407058
rect 441634 406738 441666 406974
rect 441902 406738 441986 406974
rect 442222 406738 442254 406974
rect 441634 371294 442254 406738
rect 441634 371058 441666 371294
rect 441902 371058 441986 371294
rect 442222 371058 442254 371294
rect 441634 370974 442254 371058
rect 441634 370738 441666 370974
rect 441902 370738 441986 370974
rect 442222 370738 442254 370974
rect 441634 335294 442254 370738
rect 441634 335058 441666 335294
rect 441902 335058 441986 335294
rect 442222 335058 442254 335294
rect 441634 334974 442254 335058
rect 441634 334738 441666 334974
rect 441902 334738 441986 334974
rect 442222 334738 442254 334974
rect 441634 299294 442254 334738
rect 441634 299058 441666 299294
rect 441902 299058 441986 299294
rect 442222 299058 442254 299294
rect 441634 298974 442254 299058
rect 441634 298738 441666 298974
rect 441902 298738 441986 298974
rect 442222 298738 442254 298974
rect 441634 263294 442254 298738
rect 441634 263058 441666 263294
rect 441902 263058 441986 263294
rect 442222 263058 442254 263294
rect 441634 262974 442254 263058
rect 441634 262738 441666 262974
rect 441902 262738 441986 262974
rect 442222 262738 442254 262974
rect 441634 227294 442254 262738
rect 441634 227058 441666 227294
rect 441902 227058 441986 227294
rect 442222 227058 442254 227294
rect 441634 226974 442254 227058
rect 441634 226738 441666 226974
rect 441902 226738 441986 226974
rect 442222 226738 442254 226974
rect 441634 191294 442254 226738
rect 441634 191058 441666 191294
rect 441902 191058 441986 191294
rect 442222 191058 442254 191294
rect 441634 190974 442254 191058
rect 441634 190738 441666 190974
rect 441902 190738 441986 190974
rect 442222 190738 442254 190974
rect 441634 155294 442254 190738
rect 441634 155058 441666 155294
rect 441902 155058 441986 155294
rect 442222 155058 442254 155294
rect 441634 154974 442254 155058
rect 441634 154738 441666 154974
rect 441902 154738 441986 154974
rect 442222 154738 442254 154974
rect 441634 133649 442254 154738
rect 445354 707718 445974 711590
rect 445354 707482 445386 707718
rect 445622 707482 445706 707718
rect 445942 707482 445974 707718
rect 445354 707398 445974 707482
rect 445354 707162 445386 707398
rect 445622 707162 445706 707398
rect 445942 707162 445974 707398
rect 445354 699014 445974 707162
rect 445354 698778 445386 699014
rect 445622 698778 445706 699014
rect 445942 698778 445974 699014
rect 445354 698694 445974 698778
rect 445354 698458 445386 698694
rect 445622 698458 445706 698694
rect 445942 698458 445974 698694
rect 445354 663014 445974 698458
rect 445354 662778 445386 663014
rect 445622 662778 445706 663014
rect 445942 662778 445974 663014
rect 445354 662694 445974 662778
rect 445354 662458 445386 662694
rect 445622 662458 445706 662694
rect 445942 662458 445974 662694
rect 445354 627014 445974 662458
rect 445354 626778 445386 627014
rect 445622 626778 445706 627014
rect 445942 626778 445974 627014
rect 445354 626694 445974 626778
rect 445354 626458 445386 626694
rect 445622 626458 445706 626694
rect 445942 626458 445974 626694
rect 445354 591014 445974 626458
rect 445354 590778 445386 591014
rect 445622 590778 445706 591014
rect 445942 590778 445974 591014
rect 445354 590694 445974 590778
rect 445354 590458 445386 590694
rect 445622 590458 445706 590694
rect 445942 590458 445974 590694
rect 445354 555014 445974 590458
rect 445354 554778 445386 555014
rect 445622 554778 445706 555014
rect 445942 554778 445974 555014
rect 445354 554694 445974 554778
rect 445354 554458 445386 554694
rect 445622 554458 445706 554694
rect 445942 554458 445974 554694
rect 445354 519014 445974 554458
rect 445354 518778 445386 519014
rect 445622 518778 445706 519014
rect 445942 518778 445974 519014
rect 445354 518694 445974 518778
rect 445354 518458 445386 518694
rect 445622 518458 445706 518694
rect 445942 518458 445974 518694
rect 445354 483014 445974 518458
rect 445354 482778 445386 483014
rect 445622 482778 445706 483014
rect 445942 482778 445974 483014
rect 445354 482694 445974 482778
rect 445354 482458 445386 482694
rect 445622 482458 445706 482694
rect 445942 482458 445974 482694
rect 445354 447014 445974 482458
rect 445354 446778 445386 447014
rect 445622 446778 445706 447014
rect 445942 446778 445974 447014
rect 445354 446694 445974 446778
rect 445354 446458 445386 446694
rect 445622 446458 445706 446694
rect 445942 446458 445974 446694
rect 445354 411014 445974 446458
rect 445354 410778 445386 411014
rect 445622 410778 445706 411014
rect 445942 410778 445974 411014
rect 445354 410694 445974 410778
rect 445354 410458 445386 410694
rect 445622 410458 445706 410694
rect 445942 410458 445974 410694
rect 445354 375014 445974 410458
rect 445354 374778 445386 375014
rect 445622 374778 445706 375014
rect 445942 374778 445974 375014
rect 445354 374694 445974 374778
rect 445354 374458 445386 374694
rect 445622 374458 445706 374694
rect 445942 374458 445974 374694
rect 445354 339014 445974 374458
rect 445354 338778 445386 339014
rect 445622 338778 445706 339014
rect 445942 338778 445974 339014
rect 445354 338694 445974 338778
rect 445354 338458 445386 338694
rect 445622 338458 445706 338694
rect 445942 338458 445974 338694
rect 445354 303014 445974 338458
rect 445354 302778 445386 303014
rect 445622 302778 445706 303014
rect 445942 302778 445974 303014
rect 445354 302694 445974 302778
rect 445354 302458 445386 302694
rect 445622 302458 445706 302694
rect 445942 302458 445974 302694
rect 445354 267014 445974 302458
rect 445354 266778 445386 267014
rect 445622 266778 445706 267014
rect 445942 266778 445974 267014
rect 445354 266694 445974 266778
rect 445354 266458 445386 266694
rect 445622 266458 445706 266694
rect 445942 266458 445974 266694
rect 445354 231014 445974 266458
rect 445354 230778 445386 231014
rect 445622 230778 445706 231014
rect 445942 230778 445974 231014
rect 445354 230694 445974 230778
rect 445354 230458 445386 230694
rect 445622 230458 445706 230694
rect 445942 230458 445974 230694
rect 445354 195014 445974 230458
rect 445354 194778 445386 195014
rect 445622 194778 445706 195014
rect 445942 194778 445974 195014
rect 445354 194694 445974 194778
rect 445354 194458 445386 194694
rect 445622 194458 445706 194694
rect 445942 194458 445974 194694
rect 445354 159014 445974 194458
rect 445354 158778 445386 159014
rect 445622 158778 445706 159014
rect 445942 158778 445974 159014
rect 445354 158694 445974 158778
rect 445354 158458 445386 158694
rect 445622 158458 445706 158694
rect 445942 158458 445974 158694
rect 445354 133649 445974 158458
rect 449074 708678 449694 711590
rect 449074 708442 449106 708678
rect 449342 708442 449426 708678
rect 449662 708442 449694 708678
rect 449074 708358 449694 708442
rect 449074 708122 449106 708358
rect 449342 708122 449426 708358
rect 449662 708122 449694 708358
rect 449074 666734 449694 708122
rect 449074 666498 449106 666734
rect 449342 666498 449426 666734
rect 449662 666498 449694 666734
rect 449074 666414 449694 666498
rect 449074 666178 449106 666414
rect 449342 666178 449426 666414
rect 449662 666178 449694 666414
rect 449074 630734 449694 666178
rect 449074 630498 449106 630734
rect 449342 630498 449426 630734
rect 449662 630498 449694 630734
rect 449074 630414 449694 630498
rect 449074 630178 449106 630414
rect 449342 630178 449426 630414
rect 449662 630178 449694 630414
rect 449074 594734 449694 630178
rect 449074 594498 449106 594734
rect 449342 594498 449426 594734
rect 449662 594498 449694 594734
rect 449074 594414 449694 594498
rect 449074 594178 449106 594414
rect 449342 594178 449426 594414
rect 449662 594178 449694 594414
rect 449074 558734 449694 594178
rect 449074 558498 449106 558734
rect 449342 558498 449426 558734
rect 449662 558498 449694 558734
rect 449074 558414 449694 558498
rect 449074 558178 449106 558414
rect 449342 558178 449426 558414
rect 449662 558178 449694 558414
rect 449074 522734 449694 558178
rect 449074 522498 449106 522734
rect 449342 522498 449426 522734
rect 449662 522498 449694 522734
rect 449074 522414 449694 522498
rect 449074 522178 449106 522414
rect 449342 522178 449426 522414
rect 449662 522178 449694 522414
rect 449074 486734 449694 522178
rect 449074 486498 449106 486734
rect 449342 486498 449426 486734
rect 449662 486498 449694 486734
rect 449074 486414 449694 486498
rect 449074 486178 449106 486414
rect 449342 486178 449426 486414
rect 449662 486178 449694 486414
rect 449074 450734 449694 486178
rect 449074 450498 449106 450734
rect 449342 450498 449426 450734
rect 449662 450498 449694 450734
rect 449074 450414 449694 450498
rect 449074 450178 449106 450414
rect 449342 450178 449426 450414
rect 449662 450178 449694 450414
rect 449074 414734 449694 450178
rect 449074 414498 449106 414734
rect 449342 414498 449426 414734
rect 449662 414498 449694 414734
rect 449074 414414 449694 414498
rect 449074 414178 449106 414414
rect 449342 414178 449426 414414
rect 449662 414178 449694 414414
rect 449074 378734 449694 414178
rect 449074 378498 449106 378734
rect 449342 378498 449426 378734
rect 449662 378498 449694 378734
rect 449074 378414 449694 378498
rect 449074 378178 449106 378414
rect 449342 378178 449426 378414
rect 449662 378178 449694 378414
rect 449074 342734 449694 378178
rect 449074 342498 449106 342734
rect 449342 342498 449426 342734
rect 449662 342498 449694 342734
rect 449074 342414 449694 342498
rect 449074 342178 449106 342414
rect 449342 342178 449426 342414
rect 449662 342178 449694 342414
rect 449074 306734 449694 342178
rect 449074 306498 449106 306734
rect 449342 306498 449426 306734
rect 449662 306498 449694 306734
rect 449074 306414 449694 306498
rect 449074 306178 449106 306414
rect 449342 306178 449426 306414
rect 449662 306178 449694 306414
rect 449074 270734 449694 306178
rect 449074 270498 449106 270734
rect 449342 270498 449426 270734
rect 449662 270498 449694 270734
rect 449074 270414 449694 270498
rect 449074 270178 449106 270414
rect 449342 270178 449426 270414
rect 449662 270178 449694 270414
rect 449074 234734 449694 270178
rect 449074 234498 449106 234734
rect 449342 234498 449426 234734
rect 449662 234498 449694 234734
rect 449074 234414 449694 234498
rect 449074 234178 449106 234414
rect 449342 234178 449426 234414
rect 449662 234178 449694 234414
rect 449074 198734 449694 234178
rect 449074 198498 449106 198734
rect 449342 198498 449426 198734
rect 449662 198498 449694 198734
rect 449074 198414 449694 198498
rect 449074 198178 449106 198414
rect 449342 198178 449426 198414
rect 449662 198178 449694 198414
rect 449074 162734 449694 198178
rect 449074 162498 449106 162734
rect 449342 162498 449426 162734
rect 449662 162498 449694 162734
rect 449074 162414 449694 162498
rect 449074 162178 449106 162414
rect 449342 162178 449426 162414
rect 449662 162178 449694 162414
rect 449074 133649 449694 162178
rect 452794 709638 453414 711590
rect 452794 709402 452826 709638
rect 453062 709402 453146 709638
rect 453382 709402 453414 709638
rect 452794 709318 453414 709402
rect 452794 709082 452826 709318
rect 453062 709082 453146 709318
rect 453382 709082 453414 709318
rect 452794 670454 453414 709082
rect 452794 670218 452826 670454
rect 453062 670218 453146 670454
rect 453382 670218 453414 670454
rect 452794 670134 453414 670218
rect 452794 669898 452826 670134
rect 453062 669898 453146 670134
rect 453382 669898 453414 670134
rect 452794 634454 453414 669898
rect 452794 634218 452826 634454
rect 453062 634218 453146 634454
rect 453382 634218 453414 634454
rect 452794 634134 453414 634218
rect 452794 633898 452826 634134
rect 453062 633898 453146 634134
rect 453382 633898 453414 634134
rect 452794 598454 453414 633898
rect 452794 598218 452826 598454
rect 453062 598218 453146 598454
rect 453382 598218 453414 598454
rect 452794 598134 453414 598218
rect 452794 597898 452826 598134
rect 453062 597898 453146 598134
rect 453382 597898 453414 598134
rect 452794 562454 453414 597898
rect 452794 562218 452826 562454
rect 453062 562218 453146 562454
rect 453382 562218 453414 562454
rect 452794 562134 453414 562218
rect 452794 561898 452826 562134
rect 453062 561898 453146 562134
rect 453382 561898 453414 562134
rect 452794 526454 453414 561898
rect 452794 526218 452826 526454
rect 453062 526218 453146 526454
rect 453382 526218 453414 526454
rect 452794 526134 453414 526218
rect 452794 525898 452826 526134
rect 453062 525898 453146 526134
rect 453382 525898 453414 526134
rect 452794 490454 453414 525898
rect 452794 490218 452826 490454
rect 453062 490218 453146 490454
rect 453382 490218 453414 490454
rect 452794 490134 453414 490218
rect 452794 489898 452826 490134
rect 453062 489898 453146 490134
rect 453382 489898 453414 490134
rect 452794 454454 453414 489898
rect 452794 454218 452826 454454
rect 453062 454218 453146 454454
rect 453382 454218 453414 454454
rect 452794 454134 453414 454218
rect 452794 453898 452826 454134
rect 453062 453898 453146 454134
rect 453382 453898 453414 454134
rect 452794 418454 453414 453898
rect 452794 418218 452826 418454
rect 453062 418218 453146 418454
rect 453382 418218 453414 418454
rect 452794 418134 453414 418218
rect 452794 417898 452826 418134
rect 453062 417898 453146 418134
rect 453382 417898 453414 418134
rect 452794 382454 453414 417898
rect 452794 382218 452826 382454
rect 453062 382218 453146 382454
rect 453382 382218 453414 382454
rect 452794 382134 453414 382218
rect 452794 381898 452826 382134
rect 453062 381898 453146 382134
rect 453382 381898 453414 382134
rect 452794 346454 453414 381898
rect 452794 346218 452826 346454
rect 453062 346218 453146 346454
rect 453382 346218 453414 346454
rect 452794 346134 453414 346218
rect 452794 345898 452826 346134
rect 453062 345898 453146 346134
rect 453382 345898 453414 346134
rect 452794 310454 453414 345898
rect 452794 310218 452826 310454
rect 453062 310218 453146 310454
rect 453382 310218 453414 310454
rect 452794 310134 453414 310218
rect 452794 309898 452826 310134
rect 453062 309898 453146 310134
rect 453382 309898 453414 310134
rect 452794 274454 453414 309898
rect 452794 274218 452826 274454
rect 453062 274218 453146 274454
rect 453382 274218 453414 274454
rect 452794 274134 453414 274218
rect 452794 273898 452826 274134
rect 453062 273898 453146 274134
rect 453382 273898 453414 274134
rect 452794 238454 453414 273898
rect 452794 238218 452826 238454
rect 453062 238218 453146 238454
rect 453382 238218 453414 238454
rect 452794 238134 453414 238218
rect 452794 237898 452826 238134
rect 453062 237898 453146 238134
rect 453382 237898 453414 238134
rect 452794 202454 453414 237898
rect 452794 202218 452826 202454
rect 453062 202218 453146 202454
rect 453382 202218 453414 202454
rect 452794 202134 453414 202218
rect 452794 201898 452826 202134
rect 453062 201898 453146 202134
rect 453382 201898 453414 202134
rect 452794 166454 453414 201898
rect 452794 166218 452826 166454
rect 453062 166218 453146 166454
rect 453382 166218 453414 166454
rect 452794 166134 453414 166218
rect 452794 165898 452826 166134
rect 453062 165898 453146 166134
rect 453382 165898 453414 166134
rect 420514 133586 421134 133618
rect 409354 122778 409386 123014
rect 409622 122778 409706 123014
rect 409942 122778 409974 123014
rect 409354 122694 409974 122778
rect 409354 122458 409386 122694
rect 409622 122458 409706 122694
rect 409942 122458 409974 122694
rect 409354 87014 409974 122458
rect 452794 130454 453414 165898
rect 452794 130218 452826 130454
rect 453062 130218 453146 130454
rect 453382 130218 453414 130454
rect 452794 130134 453414 130218
rect 452794 129898 452826 130134
rect 453062 129898 453146 130134
rect 453382 129898 453414 130134
rect 419568 115574 419888 115606
rect 419568 115338 419610 115574
rect 419846 115338 419888 115574
rect 419568 115254 419888 115338
rect 419568 115018 419610 115254
rect 419846 115018 419888 115254
rect 419568 114986 419888 115018
rect 450288 115574 450608 115606
rect 450288 115338 450330 115574
rect 450566 115338 450608 115574
rect 450288 115254 450608 115338
rect 450288 115018 450330 115254
rect 450566 115018 450608 115254
rect 450288 114986 450608 115018
rect 434928 111854 435248 111886
rect 434928 111618 434970 111854
rect 435206 111618 435248 111854
rect 434928 111534 435248 111618
rect 434928 111298 434970 111534
rect 435206 111298 435248 111534
rect 434928 111266 435248 111298
rect 409354 86778 409386 87014
rect 409622 86778 409706 87014
rect 409942 86778 409974 87014
rect 409354 86694 409974 86778
rect 409354 86458 409386 86694
rect 409622 86458 409706 86694
rect 409942 86458 409974 86694
rect 409091 77348 409157 77349
rect 409091 77284 409092 77348
rect 409156 77284 409157 77348
rect 409091 77283 409157 77284
rect 405634 47058 405666 47294
rect 405902 47058 405986 47294
rect 406222 47058 406254 47294
rect 405634 46974 406254 47058
rect 405634 46738 405666 46974
rect 405902 46738 405986 46974
rect 406222 46738 406254 46974
rect 405634 11294 406254 46738
rect 405634 11058 405666 11294
rect 405902 11058 405986 11294
rect 406222 11058 406254 11294
rect 405634 10974 406254 11058
rect 405634 10738 405666 10974
rect 405902 10738 405986 10974
rect 406222 10738 406254 10974
rect 405634 -2266 406254 10738
rect 409094 3773 409154 77283
rect 409354 51014 409974 86458
rect 452794 94454 453414 129898
rect 452794 94218 452826 94454
rect 453062 94218 453146 94454
rect 453382 94218 453414 94454
rect 452794 94134 453414 94218
rect 452794 93898 452826 94134
rect 453062 93898 453146 94134
rect 453382 93898 453414 94134
rect 410379 77892 410445 77893
rect 410379 77828 410380 77892
rect 410444 77828 410445 77892
rect 410379 77827 410445 77828
rect 409354 50778 409386 51014
rect 409622 50778 409706 51014
rect 409942 50778 409974 51014
rect 409354 50694 409974 50778
rect 409354 50458 409386 50694
rect 409622 50458 409706 50694
rect 409942 50458 409974 50694
rect 409354 15014 409974 50458
rect 409354 14778 409386 15014
rect 409622 14778 409706 15014
rect 409942 14778 409974 15014
rect 409354 14694 409974 14778
rect 409354 14458 409386 14694
rect 409622 14458 409706 14694
rect 409942 14458 409974 14694
rect 409091 3772 409157 3773
rect 409091 3708 409092 3772
rect 409156 3708 409157 3772
rect 409091 3707 409157 3708
rect 405634 -2502 405666 -2266
rect 405902 -2502 405986 -2266
rect 406222 -2502 406254 -2266
rect 405634 -2586 406254 -2502
rect 405634 -2822 405666 -2586
rect 405902 -2822 405986 -2586
rect 406222 -2822 406254 -2586
rect 405634 -7654 406254 -2822
rect 409354 -3226 409974 14458
rect 410382 3365 410442 77827
rect 413074 54734 413694 81159
rect 413074 54498 413106 54734
rect 413342 54498 413426 54734
rect 413662 54498 413694 54734
rect 413074 54414 413694 54498
rect 413074 54178 413106 54414
rect 413342 54178 413426 54414
rect 413662 54178 413694 54414
rect 413074 18734 413694 54178
rect 413074 18498 413106 18734
rect 413342 18498 413426 18734
rect 413662 18498 413694 18734
rect 413074 18414 413694 18498
rect 413074 18178 413106 18414
rect 413342 18178 413426 18414
rect 413662 18178 413694 18414
rect 410379 3364 410445 3365
rect 410379 3300 410380 3364
rect 410444 3300 410445 3364
rect 410379 3299 410445 3300
rect 409354 -3462 409386 -3226
rect 409622 -3462 409706 -3226
rect 409942 -3462 409974 -3226
rect 409354 -3546 409974 -3462
rect 409354 -3782 409386 -3546
rect 409622 -3782 409706 -3546
rect 409942 -3782 409974 -3546
rect 409354 -7654 409974 -3782
rect 413074 -4186 413694 18178
rect 413074 -4422 413106 -4186
rect 413342 -4422 413426 -4186
rect 413662 -4422 413694 -4186
rect 413074 -4506 413694 -4422
rect 413074 -4742 413106 -4506
rect 413342 -4742 413426 -4506
rect 413662 -4742 413694 -4506
rect 413074 -7654 413694 -4742
rect 416794 58454 417414 81159
rect 416794 58218 416826 58454
rect 417062 58218 417146 58454
rect 417382 58218 417414 58454
rect 416794 58134 417414 58218
rect 416794 57898 416826 58134
rect 417062 57898 417146 58134
rect 417382 57898 417414 58134
rect 416794 22454 417414 57898
rect 416794 22218 416826 22454
rect 417062 22218 417146 22454
rect 417382 22218 417414 22454
rect 416794 22134 417414 22218
rect 416794 21898 416826 22134
rect 417062 21898 417146 22134
rect 417382 21898 417414 22134
rect 416794 -5146 417414 21898
rect 416794 -5382 416826 -5146
rect 417062 -5382 417146 -5146
rect 417382 -5382 417414 -5146
rect 416794 -5466 417414 -5382
rect 416794 -5702 416826 -5466
rect 417062 -5702 417146 -5466
rect 417382 -5702 417414 -5466
rect 416794 -7654 417414 -5702
rect 420514 62174 421134 81159
rect 420514 61938 420546 62174
rect 420782 61938 420866 62174
rect 421102 61938 421134 62174
rect 420514 61854 421134 61938
rect 420514 61618 420546 61854
rect 420782 61618 420866 61854
rect 421102 61618 421134 61854
rect 420514 26174 421134 61618
rect 420514 25938 420546 26174
rect 420782 25938 420866 26174
rect 421102 25938 421134 26174
rect 420514 25854 421134 25938
rect 420514 25618 420546 25854
rect 420782 25618 420866 25854
rect 421102 25618 421134 25854
rect 420514 -6106 421134 25618
rect 420514 -6342 420546 -6106
rect 420782 -6342 420866 -6106
rect 421102 -6342 421134 -6106
rect 420514 -6426 421134 -6342
rect 420514 -6662 420546 -6426
rect 420782 -6662 420866 -6426
rect 421102 -6662 421134 -6426
rect 420514 -7654 421134 -6662
rect 424234 65894 424854 81159
rect 431907 78572 431973 78573
rect 431907 78570 431908 78572
rect 424234 65658 424266 65894
rect 424502 65658 424586 65894
rect 424822 65658 424854 65894
rect 424234 65574 424854 65658
rect 424234 65338 424266 65574
rect 424502 65338 424586 65574
rect 424822 65338 424854 65574
rect 424234 29894 424854 65338
rect 424234 29658 424266 29894
rect 424502 29658 424586 29894
rect 424822 29658 424854 29894
rect 424234 29574 424854 29658
rect 424234 29338 424266 29574
rect 424502 29338 424586 29574
rect 424822 29338 424854 29574
rect 424234 -7066 424854 29338
rect 431726 78510 431908 78570
rect 431726 9298 431786 78510
rect 431907 78508 431908 78510
rect 431972 78508 431973 78572
rect 431907 78507 431973 78508
rect 434194 75854 434814 79988
rect 434194 75618 434226 75854
rect 434462 75618 434546 75854
rect 434782 75618 434814 75854
rect 434194 75534 434814 75618
rect 434194 75298 434226 75534
rect 434462 75298 434546 75534
rect 434782 75298 434814 75534
rect 434194 39854 434814 75298
rect 434194 39618 434226 39854
rect 434462 39618 434546 39854
rect 434782 39618 434814 39854
rect 434194 39534 434814 39618
rect 434194 39298 434226 39534
rect 434462 39298 434546 39534
rect 434782 39298 434814 39534
rect 424234 -7302 424266 -7066
rect 424502 -7302 424586 -7066
rect 424822 -7302 424854 -7066
rect 424234 -7386 424854 -7302
rect 424234 -7622 424266 -7386
rect 424502 -7622 424586 -7386
rect 424822 -7622 424854 -7386
rect 424234 -7654 424854 -7622
rect 434194 3854 434814 39298
rect 434194 3618 434226 3854
rect 434462 3618 434546 3854
rect 434782 3618 434814 3854
rect 434194 3534 434814 3618
rect 434194 3298 434226 3534
rect 434462 3298 434546 3534
rect 434782 3298 434814 3534
rect 434194 -346 434814 3298
rect 434194 -582 434226 -346
rect 434462 -582 434546 -346
rect 434782 -582 434814 -346
rect 434194 -666 434814 -582
rect 434194 -902 434226 -666
rect 434462 -902 434546 -666
rect 434782 -902 434814 -666
rect 434194 -7654 434814 -902
rect 437914 79574 438534 81159
rect 437914 79338 437946 79574
rect 438182 79338 438266 79574
rect 438502 79338 438534 79574
rect 437914 79254 438534 79338
rect 437914 79018 437946 79254
rect 438182 79018 438266 79254
rect 438502 79018 438534 79254
rect 437914 43574 438534 79018
rect 437914 43338 437946 43574
rect 438182 43338 438266 43574
rect 438502 43338 438534 43574
rect 437914 43254 438534 43338
rect 437914 43018 437946 43254
rect 438182 43018 438266 43254
rect 438502 43018 438534 43254
rect 437914 7574 438534 43018
rect 437914 7338 437946 7574
rect 438182 7338 438266 7574
rect 438502 7338 438534 7574
rect 437914 7254 438534 7338
rect 437914 7018 437946 7254
rect 438182 7018 438266 7254
rect 438502 7018 438534 7254
rect 437914 -1306 438534 7018
rect 437914 -1542 437946 -1306
rect 438182 -1542 438266 -1306
rect 438502 -1542 438534 -1306
rect 437914 -1626 438534 -1542
rect 437914 -1862 437946 -1626
rect 438182 -1862 438266 -1626
rect 438502 -1862 438534 -1626
rect 437914 -7654 438534 -1862
rect 441634 47294 442254 81159
rect 441634 47058 441666 47294
rect 441902 47058 441986 47294
rect 442222 47058 442254 47294
rect 441634 46974 442254 47058
rect 441634 46738 441666 46974
rect 441902 46738 441986 46974
rect 442222 46738 442254 46974
rect 441634 11294 442254 46738
rect 441634 11058 441666 11294
rect 441902 11058 441986 11294
rect 442222 11058 442254 11294
rect 441634 10974 442254 11058
rect 441634 10738 441666 10974
rect 441902 10738 441986 10974
rect 442222 10738 442254 10974
rect 441634 -2266 442254 10738
rect 441634 -2502 441666 -2266
rect 441902 -2502 441986 -2266
rect 442222 -2502 442254 -2266
rect 441634 -2586 442254 -2502
rect 441634 -2822 441666 -2586
rect 441902 -2822 441986 -2586
rect 442222 -2822 442254 -2586
rect 441634 -7654 442254 -2822
rect 445354 51014 445974 81159
rect 445354 50778 445386 51014
rect 445622 50778 445706 51014
rect 445942 50778 445974 51014
rect 445354 50694 445974 50778
rect 445354 50458 445386 50694
rect 445622 50458 445706 50694
rect 445942 50458 445974 50694
rect 445354 15014 445974 50458
rect 445354 14778 445386 15014
rect 445622 14778 445706 15014
rect 445942 14778 445974 15014
rect 445354 14694 445974 14778
rect 445354 14458 445386 14694
rect 445622 14458 445706 14694
rect 445942 14458 445974 14694
rect 445354 -3226 445974 14458
rect 445354 -3462 445386 -3226
rect 445622 -3462 445706 -3226
rect 445942 -3462 445974 -3226
rect 445354 -3546 445974 -3462
rect 445354 -3782 445386 -3546
rect 445622 -3782 445706 -3546
rect 445942 -3782 445974 -3546
rect 445354 -7654 445974 -3782
rect 449074 54734 449694 81159
rect 449074 54498 449106 54734
rect 449342 54498 449426 54734
rect 449662 54498 449694 54734
rect 449074 54414 449694 54498
rect 449074 54178 449106 54414
rect 449342 54178 449426 54414
rect 449662 54178 449694 54414
rect 449074 18734 449694 54178
rect 449074 18498 449106 18734
rect 449342 18498 449426 18734
rect 449662 18498 449694 18734
rect 449074 18414 449694 18498
rect 449074 18178 449106 18414
rect 449342 18178 449426 18414
rect 449662 18178 449694 18414
rect 449074 -4186 449694 18178
rect 449074 -4422 449106 -4186
rect 449342 -4422 449426 -4186
rect 449662 -4422 449694 -4186
rect 449074 -4506 449694 -4422
rect 449074 -4742 449106 -4506
rect 449342 -4742 449426 -4506
rect 449662 -4742 449694 -4506
rect 449074 -7654 449694 -4742
rect 452794 58454 453414 93898
rect 452794 58218 452826 58454
rect 453062 58218 453146 58454
rect 453382 58218 453414 58454
rect 452794 58134 453414 58218
rect 452794 57898 452826 58134
rect 453062 57898 453146 58134
rect 453382 57898 453414 58134
rect 452794 22454 453414 57898
rect 452794 22218 452826 22454
rect 453062 22218 453146 22454
rect 453382 22218 453414 22454
rect 452794 22134 453414 22218
rect 452794 21898 452826 22134
rect 453062 21898 453146 22134
rect 453382 21898 453414 22134
rect 452794 -5146 453414 21898
rect 452794 -5382 452826 -5146
rect 453062 -5382 453146 -5146
rect 453382 -5382 453414 -5146
rect 452794 -5466 453414 -5382
rect 452794 -5702 452826 -5466
rect 453062 -5702 453146 -5466
rect 453382 -5702 453414 -5466
rect 452794 -7654 453414 -5702
rect 456514 710598 457134 711590
rect 456514 710362 456546 710598
rect 456782 710362 456866 710598
rect 457102 710362 457134 710598
rect 456514 710278 457134 710362
rect 456514 710042 456546 710278
rect 456782 710042 456866 710278
rect 457102 710042 457134 710278
rect 456514 674174 457134 710042
rect 456514 673938 456546 674174
rect 456782 673938 456866 674174
rect 457102 673938 457134 674174
rect 456514 673854 457134 673938
rect 456514 673618 456546 673854
rect 456782 673618 456866 673854
rect 457102 673618 457134 673854
rect 456514 638174 457134 673618
rect 456514 637938 456546 638174
rect 456782 637938 456866 638174
rect 457102 637938 457134 638174
rect 456514 637854 457134 637938
rect 456514 637618 456546 637854
rect 456782 637618 456866 637854
rect 457102 637618 457134 637854
rect 456514 602174 457134 637618
rect 456514 601938 456546 602174
rect 456782 601938 456866 602174
rect 457102 601938 457134 602174
rect 456514 601854 457134 601938
rect 456514 601618 456546 601854
rect 456782 601618 456866 601854
rect 457102 601618 457134 601854
rect 456514 566174 457134 601618
rect 456514 565938 456546 566174
rect 456782 565938 456866 566174
rect 457102 565938 457134 566174
rect 456514 565854 457134 565938
rect 456514 565618 456546 565854
rect 456782 565618 456866 565854
rect 457102 565618 457134 565854
rect 456514 530174 457134 565618
rect 456514 529938 456546 530174
rect 456782 529938 456866 530174
rect 457102 529938 457134 530174
rect 456514 529854 457134 529938
rect 456514 529618 456546 529854
rect 456782 529618 456866 529854
rect 457102 529618 457134 529854
rect 456514 494174 457134 529618
rect 456514 493938 456546 494174
rect 456782 493938 456866 494174
rect 457102 493938 457134 494174
rect 456514 493854 457134 493938
rect 456514 493618 456546 493854
rect 456782 493618 456866 493854
rect 457102 493618 457134 493854
rect 456514 458174 457134 493618
rect 456514 457938 456546 458174
rect 456782 457938 456866 458174
rect 457102 457938 457134 458174
rect 456514 457854 457134 457938
rect 456514 457618 456546 457854
rect 456782 457618 456866 457854
rect 457102 457618 457134 457854
rect 456514 422174 457134 457618
rect 456514 421938 456546 422174
rect 456782 421938 456866 422174
rect 457102 421938 457134 422174
rect 456514 421854 457134 421938
rect 456514 421618 456546 421854
rect 456782 421618 456866 421854
rect 457102 421618 457134 421854
rect 456514 386174 457134 421618
rect 456514 385938 456546 386174
rect 456782 385938 456866 386174
rect 457102 385938 457134 386174
rect 456514 385854 457134 385938
rect 456514 385618 456546 385854
rect 456782 385618 456866 385854
rect 457102 385618 457134 385854
rect 456514 350174 457134 385618
rect 456514 349938 456546 350174
rect 456782 349938 456866 350174
rect 457102 349938 457134 350174
rect 456514 349854 457134 349938
rect 456514 349618 456546 349854
rect 456782 349618 456866 349854
rect 457102 349618 457134 349854
rect 456514 314174 457134 349618
rect 456514 313938 456546 314174
rect 456782 313938 456866 314174
rect 457102 313938 457134 314174
rect 456514 313854 457134 313938
rect 456514 313618 456546 313854
rect 456782 313618 456866 313854
rect 457102 313618 457134 313854
rect 456514 278174 457134 313618
rect 456514 277938 456546 278174
rect 456782 277938 456866 278174
rect 457102 277938 457134 278174
rect 456514 277854 457134 277938
rect 456514 277618 456546 277854
rect 456782 277618 456866 277854
rect 457102 277618 457134 277854
rect 456514 242174 457134 277618
rect 456514 241938 456546 242174
rect 456782 241938 456866 242174
rect 457102 241938 457134 242174
rect 456514 241854 457134 241938
rect 456514 241618 456546 241854
rect 456782 241618 456866 241854
rect 457102 241618 457134 241854
rect 456514 206174 457134 241618
rect 456514 205938 456546 206174
rect 456782 205938 456866 206174
rect 457102 205938 457134 206174
rect 456514 205854 457134 205938
rect 456514 205618 456546 205854
rect 456782 205618 456866 205854
rect 457102 205618 457134 205854
rect 456514 170174 457134 205618
rect 456514 169938 456546 170174
rect 456782 169938 456866 170174
rect 457102 169938 457134 170174
rect 456514 169854 457134 169938
rect 456514 169618 456546 169854
rect 456782 169618 456866 169854
rect 457102 169618 457134 169854
rect 456514 134174 457134 169618
rect 456514 133938 456546 134174
rect 456782 133938 456866 134174
rect 457102 133938 457134 134174
rect 456514 133854 457134 133938
rect 456514 133618 456546 133854
rect 456782 133618 456866 133854
rect 457102 133618 457134 133854
rect 456514 98174 457134 133618
rect 456514 97938 456546 98174
rect 456782 97938 456866 98174
rect 457102 97938 457134 98174
rect 456514 97854 457134 97938
rect 456514 97618 456546 97854
rect 456782 97618 456866 97854
rect 457102 97618 457134 97854
rect 456514 62174 457134 97618
rect 456514 61938 456546 62174
rect 456782 61938 456866 62174
rect 457102 61938 457134 62174
rect 456514 61854 457134 61938
rect 456514 61618 456546 61854
rect 456782 61618 456866 61854
rect 457102 61618 457134 61854
rect 456514 26174 457134 61618
rect 456514 25938 456546 26174
rect 456782 25938 456866 26174
rect 457102 25938 457134 26174
rect 456514 25854 457134 25938
rect 456514 25618 456546 25854
rect 456782 25618 456866 25854
rect 457102 25618 457134 25854
rect 456514 -6106 457134 25618
rect 456514 -6342 456546 -6106
rect 456782 -6342 456866 -6106
rect 457102 -6342 457134 -6106
rect 456514 -6426 457134 -6342
rect 456514 -6662 456546 -6426
rect 456782 -6662 456866 -6426
rect 457102 -6662 457134 -6426
rect 456514 -7654 457134 -6662
rect 460234 711558 460854 711590
rect 460234 711322 460266 711558
rect 460502 711322 460586 711558
rect 460822 711322 460854 711558
rect 460234 711238 460854 711322
rect 460234 711002 460266 711238
rect 460502 711002 460586 711238
rect 460822 711002 460854 711238
rect 460234 677894 460854 711002
rect 460234 677658 460266 677894
rect 460502 677658 460586 677894
rect 460822 677658 460854 677894
rect 460234 677574 460854 677658
rect 460234 677338 460266 677574
rect 460502 677338 460586 677574
rect 460822 677338 460854 677574
rect 460234 641894 460854 677338
rect 460234 641658 460266 641894
rect 460502 641658 460586 641894
rect 460822 641658 460854 641894
rect 460234 641574 460854 641658
rect 460234 641338 460266 641574
rect 460502 641338 460586 641574
rect 460822 641338 460854 641574
rect 460234 605894 460854 641338
rect 460234 605658 460266 605894
rect 460502 605658 460586 605894
rect 460822 605658 460854 605894
rect 460234 605574 460854 605658
rect 460234 605338 460266 605574
rect 460502 605338 460586 605574
rect 460822 605338 460854 605574
rect 460234 569894 460854 605338
rect 460234 569658 460266 569894
rect 460502 569658 460586 569894
rect 460822 569658 460854 569894
rect 460234 569574 460854 569658
rect 460234 569338 460266 569574
rect 460502 569338 460586 569574
rect 460822 569338 460854 569574
rect 460234 533894 460854 569338
rect 460234 533658 460266 533894
rect 460502 533658 460586 533894
rect 460822 533658 460854 533894
rect 460234 533574 460854 533658
rect 460234 533338 460266 533574
rect 460502 533338 460586 533574
rect 460822 533338 460854 533574
rect 460234 497894 460854 533338
rect 460234 497658 460266 497894
rect 460502 497658 460586 497894
rect 460822 497658 460854 497894
rect 460234 497574 460854 497658
rect 460234 497338 460266 497574
rect 460502 497338 460586 497574
rect 460822 497338 460854 497574
rect 460234 461894 460854 497338
rect 460234 461658 460266 461894
rect 460502 461658 460586 461894
rect 460822 461658 460854 461894
rect 460234 461574 460854 461658
rect 460234 461338 460266 461574
rect 460502 461338 460586 461574
rect 460822 461338 460854 461574
rect 460234 425894 460854 461338
rect 460234 425658 460266 425894
rect 460502 425658 460586 425894
rect 460822 425658 460854 425894
rect 460234 425574 460854 425658
rect 460234 425338 460266 425574
rect 460502 425338 460586 425574
rect 460822 425338 460854 425574
rect 460234 389894 460854 425338
rect 460234 389658 460266 389894
rect 460502 389658 460586 389894
rect 460822 389658 460854 389894
rect 460234 389574 460854 389658
rect 460234 389338 460266 389574
rect 460502 389338 460586 389574
rect 460822 389338 460854 389574
rect 460234 353894 460854 389338
rect 460234 353658 460266 353894
rect 460502 353658 460586 353894
rect 460822 353658 460854 353894
rect 460234 353574 460854 353658
rect 460234 353338 460266 353574
rect 460502 353338 460586 353574
rect 460822 353338 460854 353574
rect 460234 317894 460854 353338
rect 460234 317658 460266 317894
rect 460502 317658 460586 317894
rect 460822 317658 460854 317894
rect 460234 317574 460854 317658
rect 460234 317338 460266 317574
rect 460502 317338 460586 317574
rect 460822 317338 460854 317574
rect 460234 281894 460854 317338
rect 460234 281658 460266 281894
rect 460502 281658 460586 281894
rect 460822 281658 460854 281894
rect 460234 281574 460854 281658
rect 460234 281338 460266 281574
rect 460502 281338 460586 281574
rect 460822 281338 460854 281574
rect 460234 245894 460854 281338
rect 460234 245658 460266 245894
rect 460502 245658 460586 245894
rect 460822 245658 460854 245894
rect 460234 245574 460854 245658
rect 460234 245338 460266 245574
rect 460502 245338 460586 245574
rect 460822 245338 460854 245574
rect 460234 209894 460854 245338
rect 460234 209658 460266 209894
rect 460502 209658 460586 209894
rect 460822 209658 460854 209894
rect 460234 209574 460854 209658
rect 460234 209338 460266 209574
rect 460502 209338 460586 209574
rect 460822 209338 460854 209574
rect 460234 173894 460854 209338
rect 460234 173658 460266 173894
rect 460502 173658 460586 173894
rect 460822 173658 460854 173894
rect 460234 173574 460854 173658
rect 460234 173338 460266 173574
rect 460502 173338 460586 173574
rect 460822 173338 460854 173574
rect 460234 137894 460854 173338
rect 460234 137658 460266 137894
rect 460502 137658 460586 137894
rect 460822 137658 460854 137894
rect 460234 137574 460854 137658
rect 460234 137338 460266 137574
rect 460502 137338 460586 137574
rect 460822 137338 460854 137574
rect 460234 101894 460854 137338
rect 460234 101658 460266 101894
rect 460502 101658 460586 101894
rect 460822 101658 460854 101894
rect 460234 101574 460854 101658
rect 460234 101338 460266 101574
rect 460502 101338 460586 101574
rect 460822 101338 460854 101574
rect 460234 65894 460854 101338
rect 460234 65658 460266 65894
rect 460502 65658 460586 65894
rect 460822 65658 460854 65894
rect 460234 65574 460854 65658
rect 460234 65338 460266 65574
rect 460502 65338 460586 65574
rect 460822 65338 460854 65574
rect 460234 29894 460854 65338
rect 460234 29658 460266 29894
rect 460502 29658 460586 29894
rect 460822 29658 460854 29894
rect 460234 29574 460854 29658
rect 460234 29338 460266 29574
rect 460502 29338 460586 29574
rect 460822 29338 460854 29574
rect 460234 -7066 460854 29338
rect 460234 -7302 460266 -7066
rect 460502 -7302 460586 -7066
rect 460822 -7302 460854 -7066
rect 460234 -7386 460854 -7302
rect 460234 -7622 460266 -7386
rect 460502 -7622 460586 -7386
rect 460822 -7622 460854 -7386
rect 460234 -7654 460854 -7622
rect 470194 704838 470814 711590
rect 470194 704602 470226 704838
rect 470462 704602 470546 704838
rect 470782 704602 470814 704838
rect 470194 704518 470814 704602
rect 470194 704282 470226 704518
rect 470462 704282 470546 704518
rect 470782 704282 470814 704518
rect 470194 687854 470814 704282
rect 470194 687618 470226 687854
rect 470462 687618 470546 687854
rect 470782 687618 470814 687854
rect 470194 687534 470814 687618
rect 470194 687298 470226 687534
rect 470462 687298 470546 687534
rect 470782 687298 470814 687534
rect 470194 651854 470814 687298
rect 470194 651618 470226 651854
rect 470462 651618 470546 651854
rect 470782 651618 470814 651854
rect 470194 651534 470814 651618
rect 470194 651298 470226 651534
rect 470462 651298 470546 651534
rect 470782 651298 470814 651534
rect 470194 615854 470814 651298
rect 470194 615618 470226 615854
rect 470462 615618 470546 615854
rect 470782 615618 470814 615854
rect 470194 615534 470814 615618
rect 470194 615298 470226 615534
rect 470462 615298 470546 615534
rect 470782 615298 470814 615534
rect 470194 579854 470814 615298
rect 470194 579618 470226 579854
rect 470462 579618 470546 579854
rect 470782 579618 470814 579854
rect 470194 579534 470814 579618
rect 470194 579298 470226 579534
rect 470462 579298 470546 579534
rect 470782 579298 470814 579534
rect 470194 543854 470814 579298
rect 470194 543618 470226 543854
rect 470462 543618 470546 543854
rect 470782 543618 470814 543854
rect 470194 543534 470814 543618
rect 470194 543298 470226 543534
rect 470462 543298 470546 543534
rect 470782 543298 470814 543534
rect 470194 507854 470814 543298
rect 470194 507618 470226 507854
rect 470462 507618 470546 507854
rect 470782 507618 470814 507854
rect 470194 507534 470814 507618
rect 470194 507298 470226 507534
rect 470462 507298 470546 507534
rect 470782 507298 470814 507534
rect 470194 471854 470814 507298
rect 470194 471618 470226 471854
rect 470462 471618 470546 471854
rect 470782 471618 470814 471854
rect 470194 471534 470814 471618
rect 470194 471298 470226 471534
rect 470462 471298 470546 471534
rect 470782 471298 470814 471534
rect 470194 435854 470814 471298
rect 470194 435618 470226 435854
rect 470462 435618 470546 435854
rect 470782 435618 470814 435854
rect 470194 435534 470814 435618
rect 470194 435298 470226 435534
rect 470462 435298 470546 435534
rect 470782 435298 470814 435534
rect 470194 399854 470814 435298
rect 470194 399618 470226 399854
rect 470462 399618 470546 399854
rect 470782 399618 470814 399854
rect 470194 399534 470814 399618
rect 470194 399298 470226 399534
rect 470462 399298 470546 399534
rect 470782 399298 470814 399534
rect 470194 363854 470814 399298
rect 470194 363618 470226 363854
rect 470462 363618 470546 363854
rect 470782 363618 470814 363854
rect 470194 363534 470814 363618
rect 470194 363298 470226 363534
rect 470462 363298 470546 363534
rect 470782 363298 470814 363534
rect 470194 327854 470814 363298
rect 470194 327618 470226 327854
rect 470462 327618 470546 327854
rect 470782 327618 470814 327854
rect 470194 327534 470814 327618
rect 470194 327298 470226 327534
rect 470462 327298 470546 327534
rect 470782 327298 470814 327534
rect 470194 291854 470814 327298
rect 470194 291618 470226 291854
rect 470462 291618 470546 291854
rect 470782 291618 470814 291854
rect 470194 291534 470814 291618
rect 470194 291298 470226 291534
rect 470462 291298 470546 291534
rect 470782 291298 470814 291534
rect 470194 255854 470814 291298
rect 470194 255618 470226 255854
rect 470462 255618 470546 255854
rect 470782 255618 470814 255854
rect 470194 255534 470814 255618
rect 470194 255298 470226 255534
rect 470462 255298 470546 255534
rect 470782 255298 470814 255534
rect 470194 219854 470814 255298
rect 470194 219618 470226 219854
rect 470462 219618 470546 219854
rect 470782 219618 470814 219854
rect 470194 219534 470814 219618
rect 470194 219298 470226 219534
rect 470462 219298 470546 219534
rect 470782 219298 470814 219534
rect 470194 183854 470814 219298
rect 470194 183618 470226 183854
rect 470462 183618 470546 183854
rect 470782 183618 470814 183854
rect 470194 183534 470814 183618
rect 470194 183298 470226 183534
rect 470462 183298 470546 183534
rect 470782 183298 470814 183534
rect 470194 147854 470814 183298
rect 470194 147618 470226 147854
rect 470462 147618 470546 147854
rect 470782 147618 470814 147854
rect 470194 147534 470814 147618
rect 470194 147298 470226 147534
rect 470462 147298 470546 147534
rect 470782 147298 470814 147534
rect 470194 111854 470814 147298
rect 470194 111618 470226 111854
rect 470462 111618 470546 111854
rect 470782 111618 470814 111854
rect 470194 111534 470814 111618
rect 470194 111298 470226 111534
rect 470462 111298 470546 111534
rect 470782 111298 470814 111534
rect 470194 75854 470814 111298
rect 470194 75618 470226 75854
rect 470462 75618 470546 75854
rect 470782 75618 470814 75854
rect 470194 75534 470814 75618
rect 470194 75298 470226 75534
rect 470462 75298 470546 75534
rect 470782 75298 470814 75534
rect 470194 39854 470814 75298
rect 470194 39618 470226 39854
rect 470462 39618 470546 39854
rect 470782 39618 470814 39854
rect 470194 39534 470814 39618
rect 470194 39298 470226 39534
rect 470462 39298 470546 39534
rect 470782 39298 470814 39534
rect 470194 3854 470814 39298
rect 470194 3618 470226 3854
rect 470462 3618 470546 3854
rect 470782 3618 470814 3854
rect 470194 3534 470814 3618
rect 470194 3298 470226 3534
rect 470462 3298 470546 3534
rect 470782 3298 470814 3534
rect 470194 -346 470814 3298
rect 470194 -582 470226 -346
rect 470462 -582 470546 -346
rect 470782 -582 470814 -346
rect 470194 -666 470814 -582
rect 470194 -902 470226 -666
rect 470462 -902 470546 -666
rect 470782 -902 470814 -666
rect 470194 -7654 470814 -902
rect 473914 705798 474534 711590
rect 473914 705562 473946 705798
rect 474182 705562 474266 705798
rect 474502 705562 474534 705798
rect 473914 705478 474534 705562
rect 473914 705242 473946 705478
rect 474182 705242 474266 705478
rect 474502 705242 474534 705478
rect 473914 691574 474534 705242
rect 473914 691338 473946 691574
rect 474182 691338 474266 691574
rect 474502 691338 474534 691574
rect 473914 691254 474534 691338
rect 473914 691018 473946 691254
rect 474182 691018 474266 691254
rect 474502 691018 474534 691254
rect 473914 655574 474534 691018
rect 473914 655338 473946 655574
rect 474182 655338 474266 655574
rect 474502 655338 474534 655574
rect 473914 655254 474534 655338
rect 473914 655018 473946 655254
rect 474182 655018 474266 655254
rect 474502 655018 474534 655254
rect 473914 619574 474534 655018
rect 473914 619338 473946 619574
rect 474182 619338 474266 619574
rect 474502 619338 474534 619574
rect 473914 619254 474534 619338
rect 473914 619018 473946 619254
rect 474182 619018 474266 619254
rect 474502 619018 474534 619254
rect 473914 583574 474534 619018
rect 473914 583338 473946 583574
rect 474182 583338 474266 583574
rect 474502 583338 474534 583574
rect 473914 583254 474534 583338
rect 473914 583018 473946 583254
rect 474182 583018 474266 583254
rect 474502 583018 474534 583254
rect 473914 547574 474534 583018
rect 473914 547338 473946 547574
rect 474182 547338 474266 547574
rect 474502 547338 474534 547574
rect 473914 547254 474534 547338
rect 473914 547018 473946 547254
rect 474182 547018 474266 547254
rect 474502 547018 474534 547254
rect 473914 511574 474534 547018
rect 473914 511338 473946 511574
rect 474182 511338 474266 511574
rect 474502 511338 474534 511574
rect 473914 511254 474534 511338
rect 473914 511018 473946 511254
rect 474182 511018 474266 511254
rect 474502 511018 474534 511254
rect 473914 475574 474534 511018
rect 473914 475338 473946 475574
rect 474182 475338 474266 475574
rect 474502 475338 474534 475574
rect 473914 475254 474534 475338
rect 473914 475018 473946 475254
rect 474182 475018 474266 475254
rect 474502 475018 474534 475254
rect 473914 439574 474534 475018
rect 473914 439338 473946 439574
rect 474182 439338 474266 439574
rect 474502 439338 474534 439574
rect 473914 439254 474534 439338
rect 473914 439018 473946 439254
rect 474182 439018 474266 439254
rect 474502 439018 474534 439254
rect 473914 403574 474534 439018
rect 473914 403338 473946 403574
rect 474182 403338 474266 403574
rect 474502 403338 474534 403574
rect 473914 403254 474534 403338
rect 473914 403018 473946 403254
rect 474182 403018 474266 403254
rect 474502 403018 474534 403254
rect 473914 367574 474534 403018
rect 473914 367338 473946 367574
rect 474182 367338 474266 367574
rect 474502 367338 474534 367574
rect 473914 367254 474534 367338
rect 473914 367018 473946 367254
rect 474182 367018 474266 367254
rect 474502 367018 474534 367254
rect 473914 331574 474534 367018
rect 473914 331338 473946 331574
rect 474182 331338 474266 331574
rect 474502 331338 474534 331574
rect 473914 331254 474534 331338
rect 473914 331018 473946 331254
rect 474182 331018 474266 331254
rect 474502 331018 474534 331254
rect 473914 295574 474534 331018
rect 473914 295338 473946 295574
rect 474182 295338 474266 295574
rect 474502 295338 474534 295574
rect 473914 295254 474534 295338
rect 473914 295018 473946 295254
rect 474182 295018 474266 295254
rect 474502 295018 474534 295254
rect 473914 259574 474534 295018
rect 473914 259338 473946 259574
rect 474182 259338 474266 259574
rect 474502 259338 474534 259574
rect 473914 259254 474534 259338
rect 473914 259018 473946 259254
rect 474182 259018 474266 259254
rect 474502 259018 474534 259254
rect 473914 223574 474534 259018
rect 473914 223338 473946 223574
rect 474182 223338 474266 223574
rect 474502 223338 474534 223574
rect 473914 223254 474534 223338
rect 473914 223018 473946 223254
rect 474182 223018 474266 223254
rect 474502 223018 474534 223254
rect 473914 187574 474534 223018
rect 473914 187338 473946 187574
rect 474182 187338 474266 187574
rect 474502 187338 474534 187574
rect 473914 187254 474534 187338
rect 473914 187018 473946 187254
rect 474182 187018 474266 187254
rect 474502 187018 474534 187254
rect 473914 151574 474534 187018
rect 473914 151338 473946 151574
rect 474182 151338 474266 151574
rect 474502 151338 474534 151574
rect 473914 151254 474534 151338
rect 473914 151018 473946 151254
rect 474182 151018 474266 151254
rect 474502 151018 474534 151254
rect 473914 115574 474534 151018
rect 473914 115338 473946 115574
rect 474182 115338 474266 115574
rect 474502 115338 474534 115574
rect 473914 115254 474534 115338
rect 473914 115018 473946 115254
rect 474182 115018 474266 115254
rect 474502 115018 474534 115254
rect 473914 79574 474534 115018
rect 473914 79338 473946 79574
rect 474182 79338 474266 79574
rect 474502 79338 474534 79574
rect 473914 79254 474534 79338
rect 473914 79018 473946 79254
rect 474182 79018 474266 79254
rect 474502 79018 474534 79254
rect 473914 43574 474534 79018
rect 473914 43338 473946 43574
rect 474182 43338 474266 43574
rect 474502 43338 474534 43574
rect 473914 43254 474534 43338
rect 473914 43018 473946 43254
rect 474182 43018 474266 43254
rect 474502 43018 474534 43254
rect 473914 7574 474534 43018
rect 473914 7338 473946 7574
rect 474182 7338 474266 7574
rect 474502 7338 474534 7574
rect 473914 7254 474534 7338
rect 473914 7018 473946 7254
rect 474182 7018 474266 7254
rect 474502 7018 474534 7254
rect 473914 -1306 474534 7018
rect 473914 -1542 473946 -1306
rect 474182 -1542 474266 -1306
rect 474502 -1542 474534 -1306
rect 473914 -1626 474534 -1542
rect 473914 -1862 473946 -1626
rect 474182 -1862 474266 -1626
rect 474502 -1862 474534 -1626
rect 473914 -7654 474534 -1862
rect 477634 706758 478254 711590
rect 477634 706522 477666 706758
rect 477902 706522 477986 706758
rect 478222 706522 478254 706758
rect 477634 706438 478254 706522
rect 477634 706202 477666 706438
rect 477902 706202 477986 706438
rect 478222 706202 478254 706438
rect 477634 695294 478254 706202
rect 477634 695058 477666 695294
rect 477902 695058 477986 695294
rect 478222 695058 478254 695294
rect 477634 694974 478254 695058
rect 477634 694738 477666 694974
rect 477902 694738 477986 694974
rect 478222 694738 478254 694974
rect 477634 659294 478254 694738
rect 477634 659058 477666 659294
rect 477902 659058 477986 659294
rect 478222 659058 478254 659294
rect 477634 658974 478254 659058
rect 477634 658738 477666 658974
rect 477902 658738 477986 658974
rect 478222 658738 478254 658974
rect 477634 623294 478254 658738
rect 477634 623058 477666 623294
rect 477902 623058 477986 623294
rect 478222 623058 478254 623294
rect 477634 622974 478254 623058
rect 477634 622738 477666 622974
rect 477902 622738 477986 622974
rect 478222 622738 478254 622974
rect 477634 587294 478254 622738
rect 477634 587058 477666 587294
rect 477902 587058 477986 587294
rect 478222 587058 478254 587294
rect 477634 586974 478254 587058
rect 477634 586738 477666 586974
rect 477902 586738 477986 586974
rect 478222 586738 478254 586974
rect 477634 551294 478254 586738
rect 477634 551058 477666 551294
rect 477902 551058 477986 551294
rect 478222 551058 478254 551294
rect 477634 550974 478254 551058
rect 477634 550738 477666 550974
rect 477902 550738 477986 550974
rect 478222 550738 478254 550974
rect 477634 515294 478254 550738
rect 477634 515058 477666 515294
rect 477902 515058 477986 515294
rect 478222 515058 478254 515294
rect 477634 514974 478254 515058
rect 477634 514738 477666 514974
rect 477902 514738 477986 514974
rect 478222 514738 478254 514974
rect 477634 479294 478254 514738
rect 477634 479058 477666 479294
rect 477902 479058 477986 479294
rect 478222 479058 478254 479294
rect 477634 478974 478254 479058
rect 477634 478738 477666 478974
rect 477902 478738 477986 478974
rect 478222 478738 478254 478974
rect 477634 443294 478254 478738
rect 477634 443058 477666 443294
rect 477902 443058 477986 443294
rect 478222 443058 478254 443294
rect 477634 442974 478254 443058
rect 477634 442738 477666 442974
rect 477902 442738 477986 442974
rect 478222 442738 478254 442974
rect 477634 407294 478254 442738
rect 477634 407058 477666 407294
rect 477902 407058 477986 407294
rect 478222 407058 478254 407294
rect 477634 406974 478254 407058
rect 477634 406738 477666 406974
rect 477902 406738 477986 406974
rect 478222 406738 478254 406974
rect 477634 371294 478254 406738
rect 477634 371058 477666 371294
rect 477902 371058 477986 371294
rect 478222 371058 478254 371294
rect 477634 370974 478254 371058
rect 477634 370738 477666 370974
rect 477902 370738 477986 370974
rect 478222 370738 478254 370974
rect 477634 335294 478254 370738
rect 477634 335058 477666 335294
rect 477902 335058 477986 335294
rect 478222 335058 478254 335294
rect 477634 334974 478254 335058
rect 477634 334738 477666 334974
rect 477902 334738 477986 334974
rect 478222 334738 478254 334974
rect 477634 299294 478254 334738
rect 477634 299058 477666 299294
rect 477902 299058 477986 299294
rect 478222 299058 478254 299294
rect 477634 298974 478254 299058
rect 477634 298738 477666 298974
rect 477902 298738 477986 298974
rect 478222 298738 478254 298974
rect 477634 263294 478254 298738
rect 477634 263058 477666 263294
rect 477902 263058 477986 263294
rect 478222 263058 478254 263294
rect 477634 262974 478254 263058
rect 477634 262738 477666 262974
rect 477902 262738 477986 262974
rect 478222 262738 478254 262974
rect 477634 227294 478254 262738
rect 477634 227058 477666 227294
rect 477902 227058 477986 227294
rect 478222 227058 478254 227294
rect 477634 226974 478254 227058
rect 477634 226738 477666 226974
rect 477902 226738 477986 226974
rect 478222 226738 478254 226974
rect 477634 191294 478254 226738
rect 477634 191058 477666 191294
rect 477902 191058 477986 191294
rect 478222 191058 478254 191294
rect 477634 190974 478254 191058
rect 477634 190738 477666 190974
rect 477902 190738 477986 190974
rect 478222 190738 478254 190974
rect 477634 155294 478254 190738
rect 477634 155058 477666 155294
rect 477902 155058 477986 155294
rect 478222 155058 478254 155294
rect 477634 154974 478254 155058
rect 477634 154738 477666 154974
rect 477902 154738 477986 154974
rect 478222 154738 478254 154974
rect 477634 119294 478254 154738
rect 477634 119058 477666 119294
rect 477902 119058 477986 119294
rect 478222 119058 478254 119294
rect 477634 118974 478254 119058
rect 477634 118738 477666 118974
rect 477902 118738 477986 118974
rect 478222 118738 478254 118974
rect 477634 83294 478254 118738
rect 477634 83058 477666 83294
rect 477902 83058 477986 83294
rect 478222 83058 478254 83294
rect 477634 82974 478254 83058
rect 477634 82738 477666 82974
rect 477902 82738 477986 82974
rect 478222 82738 478254 82974
rect 477634 47294 478254 82738
rect 477634 47058 477666 47294
rect 477902 47058 477986 47294
rect 478222 47058 478254 47294
rect 477634 46974 478254 47058
rect 477634 46738 477666 46974
rect 477902 46738 477986 46974
rect 478222 46738 478254 46974
rect 477634 11294 478254 46738
rect 477634 11058 477666 11294
rect 477902 11058 477986 11294
rect 478222 11058 478254 11294
rect 477634 10974 478254 11058
rect 477634 10738 477666 10974
rect 477902 10738 477986 10974
rect 478222 10738 478254 10974
rect 477634 -2266 478254 10738
rect 477634 -2502 477666 -2266
rect 477902 -2502 477986 -2266
rect 478222 -2502 478254 -2266
rect 477634 -2586 478254 -2502
rect 477634 -2822 477666 -2586
rect 477902 -2822 477986 -2586
rect 478222 -2822 478254 -2586
rect 477634 -7654 478254 -2822
rect 481354 707718 481974 711590
rect 481354 707482 481386 707718
rect 481622 707482 481706 707718
rect 481942 707482 481974 707718
rect 481354 707398 481974 707482
rect 481354 707162 481386 707398
rect 481622 707162 481706 707398
rect 481942 707162 481974 707398
rect 481354 699014 481974 707162
rect 481354 698778 481386 699014
rect 481622 698778 481706 699014
rect 481942 698778 481974 699014
rect 481354 698694 481974 698778
rect 481354 698458 481386 698694
rect 481622 698458 481706 698694
rect 481942 698458 481974 698694
rect 481354 663014 481974 698458
rect 481354 662778 481386 663014
rect 481622 662778 481706 663014
rect 481942 662778 481974 663014
rect 481354 662694 481974 662778
rect 481354 662458 481386 662694
rect 481622 662458 481706 662694
rect 481942 662458 481974 662694
rect 481354 627014 481974 662458
rect 481354 626778 481386 627014
rect 481622 626778 481706 627014
rect 481942 626778 481974 627014
rect 481354 626694 481974 626778
rect 481354 626458 481386 626694
rect 481622 626458 481706 626694
rect 481942 626458 481974 626694
rect 481354 591014 481974 626458
rect 481354 590778 481386 591014
rect 481622 590778 481706 591014
rect 481942 590778 481974 591014
rect 481354 590694 481974 590778
rect 481354 590458 481386 590694
rect 481622 590458 481706 590694
rect 481942 590458 481974 590694
rect 481354 555014 481974 590458
rect 481354 554778 481386 555014
rect 481622 554778 481706 555014
rect 481942 554778 481974 555014
rect 481354 554694 481974 554778
rect 481354 554458 481386 554694
rect 481622 554458 481706 554694
rect 481942 554458 481974 554694
rect 481354 519014 481974 554458
rect 481354 518778 481386 519014
rect 481622 518778 481706 519014
rect 481942 518778 481974 519014
rect 481354 518694 481974 518778
rect 481354 518458 481386 518694
rect 481622 518458 481706 518694
rect 481942 518458 481974 518694
rect 481354 483014 481974 518458
rect 481354 482778 481386 483014
rect 481622 482778 481706 483014
rect 481942 482778 481974 483014
rect 481354 482694 481974 482778
rect 481354 482458 481386 482694
rect 481622 482458 481706 482694
rect 481942 482458 481974 482694
rect 481354 447014 481974 482458
rect 481354 446778 481386 447014
rect 481622 446778 481706 447014
rect 481942 446778 481974 447014
rect 481354 446694 481974 446778
rect 481354 446458 481386 446694
rect 481622 446458 481706 446694
rect 481942 446458 481974 446694
rect 481354 411014 481974 446458
rect 481354 410778 481386 411014
rect 481622 410778 481706 411014
rect 481942 410778 481974 411014
rect 481354 410694 481974 410778
rect 481354 410458 481386 410694
rect 481622 410458 481706 410694
rect 481942 410458 481974 410694
rect 481354 375014 481974 410458
rect 481354 374778 481386 375014
rect 481622 374778 481706 375014
rect 481942 374778 481974 375014
rect 481354 374694 481974 374778
rect 481354 374458 481386 374694
rect 481622 374458 481706 374694
rect 481942 374458 481974 374694
rect 481354 339014 481974 374458
rect 481354 338778 481386 339014
rect 481622 338778 481706 339014
rect 481942 338778 481974 339014
rect 481354 338694 481974 338778
rect 481354 338458 481386 338694
rect 481622 338458 481706 338694
rect 481942 338458 481974 338694
rect 481354 303014 481974 338458
rect 481354 302778 481386 303014
rect 481622 302778 481706 303014
rect 481942 302778 481974 303014
rect 481354 302694 481974 302778
rect 481354 302458 481386 302694
rect 481622 302458 481706 302694
rect 481942 302458 481974 302694
rect 481354 267014 481974 302458
rect 481354 266778 481386 267014
rect 481622 266778 481706 267014
rect 481942 266778 481974 267014
rect 481354 266694 481974 266778
rect 481354 266458 481386 266694
rect 481622 266458 481706 266694
rect 481942 266458 481974 266694
rect 481354 231014 481974 266458
rect 481354 230778 481386 231014
rect 481622 230778 481706 231014
rect 481942 230778 481974 231014
rect 481354 230694 481974 230778
rect 481354 230458 481386 230694
rect 481622 230458 481706 230694
rect 481942 230458 481974 230694
rect 481354 195014 481974 230458
rect 481354 194778 481386 195014
rect 481622 194778 481706 195014
rect 481942 194778 481974 195014
rect 481354 194694 481974 194778
rect 481354 194458 481386 194694
rect 481622 194458 481706 194694
rect 481942 194458 481974 194694
rect 481354 159014 481974 194458
rect 481354 158778 481386 159014
rect 481622 158778 481706 159014
rect 481942 158778 481974 159014
rect 481354 158694 481974 158778
rect 481354 158458 481386 158694
rect 481622 158458 481706 158694
rect 481942 158458 481974 158694
rect 481354 123014 481974 158458
rect 481354 122778 481386 123014
rect 481622 122778 481706 123014
rect 481942 122778 481974 123014
rect 481354 122694 481974 122778
rect 481354 122458 481386 122694
rect 481622 122458 481706 122694
rect 481942 122458 481974 122694
rect 481354 87014 481974 122458
rect 481354 86778 481386 87014
rect 481622 86778 481706 87014
rect 481942 86778 481974 87014
rect 481354 86694 481974 86778
rect 481354 86458 481386 86694
rect 481622 86458 481706 86694
rect 481942 86458 481974 86694
rect 481354 51014 481974 86458
rect 481354 50778 481386 51014
rect 481622 50778 481706 51014
rect 481942 50778 481974 51014
rect 481354 50694 481974 50778
rect 481354 50458 481386 50694
rect 481622 50458 481706 50694
rect 481942 50458 481974 50694
rect 481354 15014 481974 50458
rect 481354 14778 481386 15014
rect 481622 14778 481706 15014
rect 481942 14778 481974 15014
rect 481354 14694 481974 14778
rect 481354 14458 481386 14694
rect 481622 14458 481706 14694
rect 481942 14458 481974 14694
rect 481354 -3226 481974 14458
rect 481354 -3462 481386 -3226
rect 481622 -3462 481706 -3226
rect 481942 -3462 481974 -3226
rect 481354 -3546 481974 -3462
rect 481354 -3782 481386 -3546
rect 481622 -3782 481706 -3546
rect 481942 -3782 481974 -3546
rect 481354 -7654 481974 -3782
rect 485074 708678 485694 711590
rect 485074 708442 485106 708678
rect 485342 708442 485426 708678
rect 485662 708442 485694 708678
rect 485074 708358 485694 708442
rect 485074 708122 485106 708358
rect 485342 708122 485426 708358
rect 485662 708122 485694 708358
rect 485074 666734 485694 708122
rect 485074 666498 485106 666734
rect 485342 666498 485426 666734
rect 485662 666498 485694 666734
rect 485074 666414 485694 666498
rect 485074 666178 485106 666414
rect 485342 666178 485426 666414
rect 485662 666178 485694 666414
rect 485074 630734 485694 666178
rect 485074 630498 485106 630734
rect 485342 630498 485426 630734
rect 485662 630498 485694 630734
rect 485074 630414 485694 630498
rect 485074 630178 485106 630414
rect 485342 630178 485426 630414
rect 485662 630178 485694 630414
rect 485074 594734 485694 630178
rect 485074 594498 485106 594734
rect 485342 594498 485426 594734
rect 485662 594498 485694 594734
rect 485074 594414 485694 594498
rect 485074 594178 485106 594414
rect 485342 594178 485426 594414
rect 485662 594178 485694 594414
rect 485074 558734 485694 594178
rect 485074 558498 485106 558734
rect 485342 558498 485426 558734
rect 485662 558498 485694 558734
rect 485074 558414 485694 558498
rect 485074 558178 485106 558414
rect 485342 558178 485426 558414
rect 485662 558178 485694 558414
rect 485074 522734 485694 558178
rect 485074 522498 485106 522734
rect 485342 522498 485426 522734
rect 485662 522498 485694 522734
rect 485074 522414 485694 522498
rect 485074 522178 485106 522414
rect 485342 522178 485426 522414
rect 485662 522178 485694 522414
rect 485074 486734 485694 522178
rect 485074 486498 485106 486734
rect 485342 486498 485426 486734
rect 485662 486498 485694 486734
rect 485074 486414 485694 486498
rect 485074 486178 485106 486414
rect 485342 486178 485426 486414
rect 485662 486178 485694 486414
rect 485074 450734 485694 486178
rect 485074 450498 485106 450734
rect 485342 450498 485426 450734
rect 485662 450498 485694 450734
rect 485074 450414 485694 450498
rect 485074 450178 485106 450414
rect 485342 450178 485426 450414
rect 485662 450178 485694 450414
rect 485074 414734 485694 450178
rect 485074 414498 485106 414734
rect 485342 414498 485426 414734
rect 485662 414498 485694 414734
rect 485074 414414 485694 414498
rect 485074 414178 485106 414414
rect 485342 414178 485426 414414
rect 485662 414178 485694 414414
rect 485074 378734 485694 414178
rect 485074 378498 485106 378734
rect 485342 378498 485426 378734
rect 485662 378498 485694 378734
rect 485074 378414 485694 378498
rect 485074 378178 485106 378414
rect 485342 378178 485426 378414
rect 485662 378178 485694 378414
rect 485074 342734 485694 378178
rect 485074 342498 485106 342734
rect 485342 342498 485426 342734
rect 485662 342498 485694 342734
rect 485074 342414 485694 342498
rect 485074 342178 485106 342414
rect 485342 342178 485426 342414
rect 485662 342178 485694 342414
rect 485074 306734 485694 342178
rect 485074 306498 485106 306734
rect 485342 306498 485426 306734
rect 485662 306498 485694 306734
rect 485074 306414 485694 306498
rect 485074 306178 485106 306414
rect 485342 306178 485426 306414
rect 485662 306178 485694 306414
rect 485074 270734 485694 306178
rect 485074 270498 485106 270734
rect 485342 270498 485426 270734
rect 485662 270498 485694 270734
rect 485074 270414 485694 270498
rect 485074 270178 485106 270414
rect 485342 270178 485426 270414
rect 485662 270178 485694 270414
rect 485074 234734 485694 270178
rect 485074 234498 485106 234734
rect 485342 234498 485426 234734
rect 485662 234498 485694 234734
rect 485074 234414 485694 234498
rect 485074 234178 485106 234414
rect 485342 234178 485426 234414
rect 485662 234178 485694 234414
rect 485074 198734 485694 234178
rect 485074 198498 485106 198734
rect 485342 198498 485426 198734
rect 485662 198498 485694 198734
rect 485074 198414 485694 198498
rect 485074 198178 485106 198414
rect 485342 198178 485426 198414
rect 485662 198178 485694 198414
rect 485074 162734 485694 198178
rect 485074 162498 485106 162734
rect 485342 162498 485426 162734
rect 485662 162498 485694 162734
rect 485074 162414 485694 162498
rect 485074 162178 485106 162414
rect 485342 162178 485426 162414
rect 485662 162178 485694 162414
rect 485074 126734 485694 162178
rect 485074 126498 485106 126734
rect 485342 126498 485426 126734
rect 485662 126498 485694 126734
rect 485074 126414 485694 126498
rect 485074 126178 485106 126414
rect 485342 126178 485426 126414
rect 485662 126178 485694 126414
rect 485074 90734 485694 126178
rect 485074 90498 485106 90734
rect 485342 90498 485426 90734
rect 485662 90498 485694 90734
rect 485074 90414 485694 90498
rect 485074 90178 485106 90414
rect 485342 90178 485426 90414
rect 485662 90178 485694 90414
rect 485074 54734 485694 90178
rect 485074 54498 485106 54734
rect 485342 54498 485426 54734
rect 485662 54498 485694 54734
rect 485074 54414 485694 54498
rect 485074 54178 485106 54414
rect 485342 54178 485426 54414
rect 485662 54178 485694 54414
rect 485074 18734 485694 54178
rect 485074 18498 485106 18734
rect 485342 18498 485426 18734
rect 485662 18498 485694 18734
rect 485074 18414 485694 18498
rect 485074 18178 485106 18414
rect 485342 18178 485426 18414
rect 485662 18178 485694 18414
rect 485074 -4186 485694 18178
rect 485074 -4422 485106 -4186
rect 485342 -4422 485426 -4186
rect 485662 -4422 485694 -4186
rect 485074 -4506 485694 -4422
rect 485074 -4742 485106 -4506
rect 485342 -4742 485426 -4506
rect 485662 -4742 485694 -4506
rect 485074 -7654 485694 -4742
rect 488794 709638 489414 711590
rect 488794 709402 488826 709638
rect 489062 709402 489146 709638
rect 489382 709402 489414 709638
rect 488794 709318 489414 709402
rect 488794 709082 488826 709318
rect 489062 709082 489146 709318
rect 489382 709082 489414 709318
rect 488794 670454 489414 709082
rect 488794 670218 488826 670454
rect 489062 670218 489146 670454
rect 489382 670218 489414 670454
rect 488794 670134 489414 670218
rect 488794 669898 488826 670134
rect 489062 669898 489146 670134
rect 489382 669898 489414 670134
rect 488794 634454 489414 669898
rect 488794 634218 488826 634454
rect 489062 634218 489146 634454
rect 489382 634218 489414 634454
rect 488794 634134 489414 634218
rect 488794 633898 488826 634134
rect 489062 633898 489146 634134
rect 489382 633898 489414 634134
rect 488794 598454 489414 633898
rect 488794 598218 488826 598454
rect 489062 598218 489146 598454
rect 489382 598218 489414 598454
rect 488794 598134 489414 598218
rect 488794 597898 488826 598134
rect 489062 597898 489146 598134
rect 489382 597898 489414 598134
rect 488794 562454 489414 597898
rect 488794 562218 488826 562454
rect 489062 562218 489146 562454
rect 489382 562218 489414 562454
rect 488794 562134 489414 562218
rect 488794 561898 488826 562134
rect 489062 561898 489146 562134
rect 489382 561898 489414 562134
rect 488794 526454 489414 561898
rect 488794 526218 488826 526454
rect 489062 526218 489146 526454
rect 489382 526218 489414 526454
rect 488794 526134 489414 526218
rect 488794 525898 488826 526134
rect 489062 525898 489146 526134
rect 489382 525898 489414 526134
rect 488794 490454 489414 525898
rect 488794 490218 488826 490454
rect 489062 490218 489146 490454
rect 489382 490218 489414 490454
rect 488794 490134 489414 490218
rect 488794 489898 488826 490134
rect 489062 489898 489146 490134
rect 489382 489898 489414 490134
rect 488794 454454 489414 489898
rect 488794 454218 488826 454454
rect 489062 454218 489146 454454
rect 489382 454218 489414 454454
rect 488794 454134 489414 454218
rect 488794 453898 488826 454134
rect 489062 453898 489146 454134
rect 489382 453898 489414 454134
rect 488794 418454 489414 453898
rect 488794 418218 488826 418454
rect 489062 418218 489146 418454
rect 489382 418218 489414 418454
rect 488794 418134 489414 418218
rect 488794 417898 488826 418134
rect 489062 417898 489146 418134
rect 489382 417898 489414 418134
rect 488794 382454 489414 417898
rect 488794 382218 488826 382454
rect 489062 382218 489146 382454
rect 489382 382218 489414 382454
rect 488794 382134 489414 382218
rect 488794 381898 488826 382134
rect 489062 381898 489146 382134
rect 489382 381898 489414 382134
rect 488794 346454 489414 381898
rect 488794 346218 488826 346454
rect 489062 346218 489146 346454
rect 489382 346218 489414 346454
rect 488794 346134 489414 346218
rect 488794 345898 488826 346134
rect 489062 345898 489146 346134
rect 489382 345898 489414 346134
rect 488794 310454 489414 345898
rect 488794 310218 488826 310454
rect 489062 310218 489146 310454
rect 489382 310218 489414 310454
rect 488794 310134 489414 310218
rect 488794 309898 488826 310134
rect 489062 309898 489146 310134
rect 489382 309898 489414 310134
rect 488794 274454 489414 309898
rect 488794 274218 488826 274454
rect 489062 274218 489146 274454
rect 489382 274218 489414 274454
rect 488794 274134 489414 274218
rect 488794 273898 488826 274134
rect 489062 273898 489146 274134
rect 489382 273898 489414 274134
rect 488794 238454 489414 273898
rect 488794 238218 488826 238454
rect 489062 238218 489146 238454
rect 489382 238218 489414 238454
rect 488794 238134 489414 238218
rect 488794 237898 488826 238134
rect 489062 237898 489146 238134
rect 489382 237898 489414 238134
rect 488794 202454 489414 237898
rect 488794 202218 488826 202454
rect 489062 202218 489146 202454
rect 489382 202218 489414 202454
rect 488794 202134 489414 202218
rect 488794 201898 488826 202134
rect 489062 201898 489146 202134
rect 489382 201898 489414 202134
rect 488794 166454 489414 201898
rect 488794 166218 488826 166454
rect 489062 166218 489146 166454
rect 489382 166218 489414 166454
rect 488794 166134 489414 166218
rect 488794 165898 488826 166134
rect 489062 165898 489146 166134
rect 489382 165898 489414 166134
rect 488794 130454 489414 165898
rect 488794 130218 488826 130454
rect 489062 130218 489146 130454
rect 489382 130218 489414 130454
rect 488794 130134 489414 130218
rect 488794 129898 488826 130134
rect 489062 129898 489146 130134
rect 489382 129898 489414 130134
rect 488794 94454 489414 129898
rect 488794 94218 488826 94454
rect 489062 94218 489146 94454
rect 489382 94218 489414 94454
rect 488794 94134 489414 94218
rect 488794 93898 488826 94134
rect 489062 93898 489146 94134
rect 489382 93898 489414 94134
rect 488794 58454 489414 93898
rect 488794 58218 488826 58454
rect 489062 58218 489146 58454
rect 489382 58218 489414 58454
rect 488794 58134 489414 58218
rect 488794 57898 488826 58134
rect 489062 57898 489146 58134
rect 489382 57898 489414 58134
rect 488794 22454 489414 57898
rect 488794 22218 488826 22454
rect 489062 22218 489146 22454
rect 489382 22218 489414 22454
rect 488794 22134 489414 22218
rect 488794 21898 488826 22134
rect 489062 21898 489146 22134
rect 489382 21898 489414 22134
rect 488794 -5146 489414 21898
rect 488794 -5382 488826 -5146
rect 489062 -5382 489146 -5146
rect 489382 -5382 489414 -5146
rect 488794 -5466 489414 -5382
rect 488794 -5702 488826 -5466
rect 489062 -5702 489146 -5466
rect 489382 -5702 489414 -5466
rect 488794 -7654 489414 -5702
rect 492514 710598 493134 711590
rect 492514 710362 492546 710598
rect 492782 710362 492866 710598
rect 493102 710362 493134 710598
rect 492514 710278 493134 710362
rect 492514 710042 492546 710278
rect 492782 710042 492866 710278
rect 493102 710042 493134 710278
rect 492514 674174 493134 710042
rect 492514 673938 492546 674174
rect 492782 673938 492866 674174
rect 493102 673938 493134 674174
rect 492514 673854 493134 673938
rect 492514 673618 492546 673854
rect 492782 673618 492866 673854
rect 493102 673618 493134 673854
rect 492514 638174 493134 673618
rect 492514 637938 492546 638174
rect 492782 637938 492866 638174
rect 493102 637938 493134 638174
rect 492514 637854 493134 637938
rect 492514 637618 492546 637854
rect 492782 637618 492866 637854
rect 493102 637618 493134 637854
rect 492514 602174 493134 637618
rect 492514 601938 492546 602174
rect 492782 601938 492866 602174
rect 493102 601938 493134 602174
rect 492514 601854 493134 601938
rect 492514 601618 492546 601854
rect 492782 601618 492866 601854
rect 493102 601618 493134 601854
rect 492514 566174 493134 601618
rect 492514 565938 492546 566174
rect 492782 565938 492866 566174
rect 493102 565938 493134 566174
rect 492514 565854 493134 565938
rect 492514 565618 492546 565854
rect 492782 565618 492866 565854
rect 493102 565618 493134 565854
rect 492514 530174 493134 565618
rect 492514 529938 492546 530174
rect 492782 529938 492866 530174
rect 493102 529938 493134 530174
rect 492514 529854 493134 529938
rect 492514 529618 492546 529854
rect 492782 529618 492866 529854
rect 493102 529618 493134 529854
rect 492514 494174 493134 529618
rect 492514 493938 492546 494174
rect 492782 493938 492866 494174
rect 493102 493938 493134 494174
rect 492514 493854 493134 493938
rect 492514 493618 492546 493854
rect 492782 493618 492866 493854
rect 493102 493618 493134 493854
rect 492514 458174 493134 493618
rect 492514 457938 492546 458174
rect 492782 457938 492866 458174
rect 493102 457938 493134 458174
rect 492514 457854 493134 457938
rect 492514 457618 492546 457854
rect 492782 457618 492866 457854
rect 493102 457618 493134 457854
rect 492514 422174 493134 457618
rect 492514 421938 492546 422174
rect 492782 421938 492866 422174
rect 493102 421938 493134 422174
rect 492514 421854 493134 421938
rect 492514 421618 492546 421854
rect 492782 421618 492866 421854
rect 493102 421618 493134 421854
rect 492514 386174 493134 421618
rect 492514 385938 492546 386174
rect 492782 385938 492866 386174
rect 493102 385938 493134 386174
rect 492514 385854 493134 385938
rect 492514 385618 492546 385854
rect 492782 385618 492866 385854
rect 493102 385618 493134 385854
rect 492514 350174 493134 385618
rect 492514 349938 492546 350174
rect 492782 349938 492866 350174
rect 493102 349938 493134 350174
rect 492514 349854 493134 349938
rect 492514 349618 492546 349854
rect 492782 349618 492866 349854
rect 493102 349618 493134 349854
rect 492514 314174 493134 349618
rect 492514 313938 492546 314174
rect 492782 313938 492866 314174
rect 493102 313938 493134 314174
rect 492514 313854 493134 313938
rect 492514 313618 492546 313854
rect 492782 313618 492866 313854
rect 493102 313618 493134 313854
rect 492514 278174 493134 313618
rect 492514 277938 492546 278174
rect 492782 277938 492866 278174
rect 493102 277938 493134 278174
rect 492514 277854 493134 277938
rect 492514 277618 492546 277854
rect 492782 277618 492866 277854
rect 493102 277618 493134 277854
rect 492514 242174 493134 277618
rect 492514 241938 492546 242174
rect 492782 241938 492866 242174
rect 493102 241938 493134 242174
rect 492514 241854 493134 241938
rect 492514 241618 492546 241854
rect 492782 241618 492866 241854
rect 493102 241618 493134 241854
rect 492514 206174 493134 241618
rect 492514 205938 492546 206174
rect 492782 205938 492866 206174
rect 493102 205938 493134 206174
rect 492514 205854 493134 205938
rect 492514 205618 492546 205854
rect 492782 205618 492866 205854
rect 493102 205618 493134 205854
rect 492514 170174 493134 205618
rect 492514 169938 492546 170174
rect 492782 169938 492866 170174
rect 493102 169938 493134 170174
rect 492514 169854 493134 169938
rect 492514 169618 492546 169854
rect 492782 169618 492866 169854
rect 493102 169618 493134 169854
rect 492514 134174 493134 169618
rect 492514 133938 492546 134174
rect 492782 133938 492866 134174
rect 493102 133938 493134 134174
rect 492514 133854 493134 133938
rect 492514 133618 492546 133854
rect 492782 133618 492866 133854
rect 493102 133618 493134 133854
rect 492514 98174 493134 133618
rect 492514 97938 492546 98174
rect 492782 97938 492866 98174
rect 493102 97938 493134 98174
rect 492514 97854 493134 97938
rect 492514 97618 492546 97854
rect 492782 97618 492866 97854
rect 493102 97618 493134 97854
rect 492514 62174 493134 97618
rect 492514 61938 492546 62174
rect 492782 61938 492866 62174
rect 493102 61938 493134 62174
rect 492514 61854 493134 61938
rect 492514 61618 492546 61854
rect 492782 61618 492866 61854
rect 493102 61618 493134 61854
rect 492514 26174 493134 61618
rect 492514 25938 492546 26174
rect 492782 25938 492866 26174
rect 493102 25938 493134 26174
rect 492514 25854 493134 25938
rect 492514 25618 492546 25854
rect 492782 25618 492866 25854
rect 493102 25618 493134 25854
rect 492514 -6106 493134 25618
rect 492514 -6342 492546 -6106
rect 492782 -6342 492866 -6106
rect 493102 -6342 493134 -6106
rect 492514 -6426 493134 -6342
rect 492514 -6662 492546 -6426
rect 492782 -6662 492866 -6426
rect 493102 -6662 493134 -6426
rect 492514 -7654 493134 -6662
rect 496234 711558 496854 711590
rect 496234 711322 496266 711558
rect 496502 711322 496586 711558
rect 496822 711322 496854 711558
rect 496234 711238 496854 711322
rect 496234 711002 496266 711238
rect 496502 711002 496586 711238
rect 496822 711002 496854 711238
rect 496234 677894 496854 711002
rect 496234 677658 496266 677894
rect 496502 677658 496586 677894
rect 496822 677658 496854 677894
rect 496234 677574 496854 677658
rect 496234 677338 496266 677574
rect 496502 677338 496586 677574
rect 496822 677338 496854 677574
rect 496234 641894 496854 677338
rect 496234 641658 496266 641894
rect 496502 641658 496586 641894
rect 496822 641658 496854 641894
rect 496234 641574 496854 641658
rect 496234 641338 496266 641574
rect 496502 641338 496586 641574
rect 496822 641338 496854 641574
rect 496234 605894 496854 641338
rect 496234 605658 496266 605894
rect 496502 605658 496586 605894
rect 496822 605658 496854 605894
rect 496234 605574 496854 605658
rect 496234 605338 496266 605574
rect 496502 605338 496586 605574
rect 496822 605338 496854 605574
rect 496234 569894 496854 605338
rect 496234 569658 496266 569894
rect 496502 569658 496586 569894
rect 496822 569658 496854 569894
rect 496234 569574 496854 569658
rect 496234 569338 496266 569574
rect 496502 569338 496586 569574
rect 496822 569338 496854 569574
rect 496234 533894 496854 569338
rect 496234 533658 496266 533894
rect 496502 533658 496586 533894
rect 496822 533658 496854 533894
rect 496234 533574 496854 533658
rect 496234 533338 496266 533574
rect 496502 533338 496586 533574
rect 496822 533338 496854 533574
rect 496234 497894 496854 533338
rect 496234 497658 496266 497894
rect 496502 497658 496586 497894
rect 496822 497658 496854 497894
rect 496234 497574 496854 497658
rect 496234 497338 496266 497574
rect 496502 497338 496586 497574
rect 496822 497338 496854 497574
rect 496234 461894 496854 497338
rect 496234 461658 496266 461894
rect 496502 461658 496586 461894
rect 496822 461658 496854 461894
rect 496234 461574 496854 461658
rect 496234 461338 496266 461574
rect 496502 461338 496586 461574
rect 496822 461338 496854 461574
rect 496234 425894 496854 461338
rect 496234 425658 496266 425894
rect 496502 425658 496586 425894
rect 496822 425658 496854 425894
rect 496234 425574 496854 425658
rect 496234 425338 496266 425574
rect 496502 425338 496586 425574
rect 496822 425338 496854 425574
rect 496234 389894 496854 425338
rect 496234 389658 496266 389894
rect 496502 389658 496586 389894
rect 496822 389658 496854 389894
rect 496234 389574 496854 389658
rect 496234 389338 496266 389574
rect 496502 389338 496586 389574
rect 496822 389338 496854 389574
rect 496234 353894 496854 389338
rect 496234 353658 496266 353894
rect 496502 353658 496586 353894
rect 496822 353658 496854 353894
rect 496234 353574 496854 353658
rect 496234 353338 496266 353574
rect 496502 353338 496586 353574
rect 496822 353338 496854 353574
rect 496234 317894 496854 353338
rect 496234 317658 496266 317894
rect 496502 317658 496586 317894
rect 496822 317658 496854 317894
rect 496234 317574 496854 317658
rect 496234 317338 496266 317574
rect 496502 317338 496586 317574
rect 496822 317338 496854 317574
rect 496234 281894 496854 317338
rect 496234 281658 496266 281894
rect 496502 281658 496586 281894
rect 496822 281658 496854 281894
rect 496234 281574 496854 281658
rect 496234 281338 496266 281574
rect 496502 281338 496586 281574
rect 496822 281338 496854 281574
rect 496234 245894 496854 281338
rect 496234 245658 496266 245894
rect 496502 245658 496586 245894
rect 496822 245658 496854 245894
rect 496234 245574 496854 245658
rect 496234 245338 496266 245574
rect 496502 245338 496586 245574
rect 496822 245338 496854 245574
rect 496234 209894 496854 245338
rect 496234 209658 496266 209894
rect 496502 209658 496586 209894
rect 496822 209658 496854 209894
rect 496234 209574 496854 209658
rect 496234 209338 496266 209574
rect 496502 209338 496586 209574
rect 496822 209338 496854 209574
rect 496234 173894 496854 209338
rect 496234 173658 496266 173894
rect 496502 173658 496586 173894
rect 496822 173658 496854 173894
rect 496234 173574 496854 173658
rect 496234 173338 496266 173574
rect 496502 173338 496586 173574
rect 496822 173338 496854 173574
rect 496234 137894 496854 173338
rect 496234 137658 496266 137894
rect 496502 137658 496586 137894
rect 496822 137658 496854 137894
rect 496234 137574 496854 137658
rect 496234 137338 496266 137574
rect 496502 137338 496586 137574
rect 496822 137338 496854 137574
rect 496234 101894 496854 137338
rect 496234 101658 496266 101894
rect 496502 101658 496586 101894
rect 496822 101658 496854 101894
rect 496234 101574 496854 101658
rect 496234 101338 496266 101574
rect 496502 101338 496586 101574
rect 496822 101338 496854 101574
rect 496234 65894 496854 101338
rect 496234 65658 496266 65894
rect 496502 65658 496586 65894
rect 496822 65658 496854 65894
rect 496234 65574 496854 65658
rect 496234 65338 496266 65574
rect 496502 65338 496586 65574
rect 496822 65338 496854 65574
rect 496234 29894 496854 65338
rect 496234 29658 496266 29894
rect 496502 29658 496586 29894
rect 496822 29658 496854 29894
rect 496234 29574 496854 29658
rect 496234 29338 496266 29574
rect 496502 29338 496586 29574
rect 496822 29338 496854 29574
rect 496234 -7066 496854 29338
rect 496234 -7302 496266 -7066
rect 496502 -7302 496586 -7066
rect 496822 -7302 496854 -7066
rect 496234 -7386 496854 -7302
rect 496234 -7622 496266 -7386
rect 496502 -7622 496586 -7386
rect 496822 -7622 496854 -7386
rect 496234 -7654 496854 -7622
rect 506194 704838 506814 711590
rect 506194 704602 506226 704838
rect 506462 704602 506546 704838
rect 506782 704602 506814 704838
rect 506194 704518 506814 704602
rect 506194 704282 506226 704518
rect 506462 704282 506546 704518
rect 506782 704282 506814 704518
rect 506194 687854 506814 704282
rect 506194 687618 506226 687854
rect 506462 687618 506546 687854
rect 506782 687618 506814 687854
rect 506194 687534 506814 687618
rect 506194 687298 506226 687534
rect 506462 687298 506546 687534
rect 506782 687298 506814 687534
rect 506194 651854 506814 687298
rect 506194 651618 506226 651854
rect 506462 651618 506546 651854
rect 506782 651618 506814 651854
rect 506194 651534 506814 651618
rect 506194 651298 506226 651534
rect 506462 651298 506546 651534
rect 506782 651298 506814 651534
rect 506194 615854 506814 651298
rect 506194 615618 506226 615854
rect 506462 615618 506546 615854
rect 506782 615618 506814 615854
rect 506194 615534 506814 615618
rect 506194 615298 506226 615534
rect 506462 615298 506546 615534
rect 506782 615298 506814 615534
rect 506194 579854 506814 615298
rect 506194 579618 506226 579854
rect 506462 579618 506546 579854
rect 506782 579618 506814 579854
rect 506194 579534 506814 579618
rect 506194 579298 506226 579534
rect 506462 579298 506546 579534
rect 506782 579298 506814 579534
rect 506194 543854 506814 579298
rect 506194 543618 506226 543854
rect 506462 543618 506546 543854
rect 506782 543618 506814 543854
rect 506194 543534 506814 543618
rect 506194 543298 506226 543534
rect 506462 543298 506546 543534
rect 506782 543298 506814 543534
rect 506194 507854 506814 543298
rect 506194 507618 506226 507854
rect 506462 507618 506546 507854
rect 506782 507618 506814 507854
rect 506194 507534 506814 507618
rect 506194 507298 506226 507534
rect 506462 507298 506546 507534
rect 506782 507298 506814 507534
rect 506194 471854 506814 507298
rect 506194 471618 506226 471854
rect 506462 471618 506546 471854
rect 506782 471618 506814 471854
rect 506194 471534 506814 471618
rect 506194 471298 506226 471534
rect 506462 471298 506546 471534
rect 506782 471298 506814 471534
rect 506194 435854 506814 471298
rect 506194 435618 506226 435854
rect 506462 435618 506546 435854
rect 506782 435618 506814 435854
rect 506194 435534 506814 435618
rect 506194 435298 506226 435534
rect 506462 435298 506546 435534
rect 506782 435298 506814 435534
rect 506194 399854 506814 435298
rect 506194 399618 506226 399854
rect 506462 399618 506546 399854
rect 506782 399618 506814 399854
rect 506194 399534 506814 399618
rect 506194 399298 506226 399534
rect 506462 399298 506546 399534
rect 506782 399298 506814 399534
rect 506194 363854 506814 399298
rect 506194 363618 506226 363854
rect 506462 363618 506546 363854
rect 506782 363618 506814 363854
rect 506194 363534 506814 363618
rect 506194 363298 506226 363534
rect 506462 363298 506546 363534
rect 506782 363298 506814 363534
rect 506194 327854 506814 363298
rect 506194 327618 506226 327854
rect 506462 327618 506546 327854
rect 506782 327618 506814 327854
rect 506194 327534 506814 327618
rect 506194 327298 506226 327534
rect 506462 327298 506546 327534
rect 506782 327298 506814 327534
rect 506194 291854 506814 327298
rect 506194 291618 506226 291854
rect 506462 291618 506546 291854
rect 506782 291618 506814 291854
rect 506194 291534 506814 291618
rect 506194 291298 506226 291534
rect 506462 291298 506546 291534
rect 506782 291298 506814 291534
rect 506194 255854 506814 291298
rect 506194 255618 506226 255854
rect 506462 255618 506546 255854
rect 506782 255618 506814 255854
rect 506194 255534 506814 255618
rect 506194 255298 506226 255534
rect 506462 255298 506546 255534
rect 506782 255298 506814 255534
rect 506194 219854 506814 255298
rect 506194 219618 506226 219854
rect 506462 219618 506546 219854
rect 506782 219618 506814 219854
rect 506194 219534 506814 219618
rect 506194 219298 506226 219534
rect 506462 219298 506546 219534
rect 506782 219298 506814 219534
rect 506194 183854 506814 219298
rect 506194 183618 506226 183854
rect 506462 183618 506546 183854
rect 506782 183618 506814 183854
rect 506194 183534 506814 183618
rect 506194 183298 506226 183534
rect 506462 183298 506546 183534
rect 506782 183298 506814 183534
rect 506194 147854 506814 183298
rect 506194 147618 506226 147854
rect 506462 147618 506546 147854
rect 506782 147618 506814 147854
rect 506194 147534 506814 147618
rect 506194 147298 506226 147534
rect 506462 147298 506546 147534
rect 506782 147298 506814 147534
rect 506194 111854 506814 147298
rect 506194 111618 506226 111854
rect 506462 111618 506546 111854
rect 506782 111618 506814 111854
rect 506194 111534 506814 111618
rect 506194 111298 506226 111534
rect 506462 111298 506546 111534
rect 506782 111298 506814 111534
rect 506194 75854 506814 111298
rect 506194 75618 506226 75854
rect 506462 75618 506546 75854
rect 506782 75618 506814 75854
rect 506194 75534 506814 75618
rect 506194 75298 506226 75534
rect 506462 75298 506546 75534
rect 506782 75298 506814 75534
rect 506194 39854 506814 75298
rect 506194 39618 506226 39854
rect 506462 39618 506546 39854
rect 506782 39618 506814 39854
rect 506194 39534 506814 39618
rect 506194 39298 506226 39534
rect 506462 39298 506546 39534
rect 506782 39298 506814 39534
rect 506194 3854 506814 39298
rect 506194 3618 506226 3854
rect 506462 3618 506546 3854
rect 506782 3618 506814 3854
rect 506194 3534 506814 3618
rect 506194 3298 506226 3534
rect 506462 3298 506546 3534
rect 506782 3298 506814 3534
rect 506194 -346 506814 3298
rect 506194 -582 506226 -346
rect 506462 -582 506546 -346
rect 506782 -582 506814 -346
rect 506194 -666 506814 -582
rect 506194 -902 506226 -666
rect 506462 -902 506546 -666
rect 506782 -902 506814 -666
rect 506194 -7654 506814 -902
rect 509914 705798 510534 711590
rect 509914 705562 509946 705798
rect 510182 705562 510266 705798
rect 510502 705562 510534 705798
rect 509914 705478 510534 705562
rect 509914 705242 509946 705478
rect 510182 705242 510266 705478
rect 510502 705242 510534 705478
rect 509914 691574 510534 705242
rect 509914 691338 509946 691574
rect 510182 691338 510266 691574
rect 510502 691338 510534 691574
rect 509914 691254 510534 691338
rect 509914 691018 509946 691254
rect 510182 691018 510266 691254
rect 510502 691018 510534 691254
rect 509914 655574 510534 691018
rect 509914 655338 509946 655574
rect 510182 655338 510266 655574
rect 510502 655338 510534 655574
rect 509914 655254 510534 655338
rect 509914 655018 509946 655254
rect 510182 655018 510266 655254
rect 510502 655018 510534 655254
rect 509914 619574 510534 655018
rect 509914 619338 509946 619574
rect 510182 619338 510266 619574
rect 510502 619338 510534 619574
rect 509914 619254 510534 619338
rect 509914 619018 509946 619254
rect 510182 619018 510266 619254
rect 510502 619018 510534 619254
rect 509914 583574 510534 619018
rect 509914 583338 509946 583574
rect 510182 583338 510266 583574
rect 510502 583338 510534 583574
rect 509914 583254 510534 583338
rect 509914 583018 509946 583254
rect 510182 583018 510266 583254
rect 510502 583018 510534 583254
rect 509914 547574 510534 583018
rect 509914 547338 509946 547574
rect 510182 547338 510266 547574
rect 510502 547338 510534 547574
rect 509914 547254 510534 547338
rect 509914 547018 509946 547254
rect 510182 547018 510266 547254
rect 510502 547018 510534 547254
rect 509914 511574 510534 547018
rect 509914 511338 509946 511574
rect 510182 511338 510266 511574
rect 510502 511338 510534 511574
rect 509914 511254 510534 511338
rect 509914 511018 509946 511254
rect 510182 511018 510266 511254
rect 510502 511018 510534 511254
rect 509914 475574 510534 511018
rect 509914 475338 509946 475574
rect 510182 475338 510266 475574
rect 510502 475338 510534 475574
rect 509914 475254 510534 475338
rect 509914 475018 509946 475254
rect 510182 475018 510266 475254
rect 510502 475018 510534 475254
rect 509914 439574 510534 475018
rect 509914 439338 509946 439574
rect 510182 439338 510266 439574
rect 510502 439338 510534 439574
rect 509914 439254 510534 439338
rect 509914 439018 509946 439254
rect 510182 439018 510266 439254
rect 510502 439018 510534 439254
rect 509914 403574 510534 439018
rect 509914 403338 509946 403574
rect 510182 403338 510266 403574
rect 510502 403338 510534 403574
rect 509914 403254 510534 403338
rect 509914 403018 509946 403254
rect 510182 403018 510266 403254
rect 510502 403018 510534 403254
rect 509914 367574 510534 403018
rect 509914 367338 509946 367574
rect 510182 367338 510266 367574
rect 510502 367338 510534 367574
rect 509914 367254 510534 367338
rect 509914 367018 509946 367254
rect 510182 367018 510266 367254
rect 510502 367018 510534 367254
rect 509914 331574 510534 367018
rect 509914 331338 509946 331574
rect 510182 331338 510266 331574
rect 510502 331338 510534 331574
rect 509914 331254 510534 331338
rect 509914 331018 509946 331254
rect 510182 331018 510266 331254
rect 510502 331018 510534 331254
rect 509914 295574 510534 331018
rect 509914 295338 509946 295574
rect 510182 295338 510266 295574
rect 510502 295338 510534 295574
rect 509914 295254 510534 295338
rect 509914 295018 509946 295254
rect 510182 295018 510266 295254
rect 510502 295018 510534 295254
rect 509914 259574 510534 295018
rect 509914 259338 509946 259574
rect 510182 259338 510266 259574
rect 510502 259338 510534 259574
rect 509914 259254 510534 259338
rect 509914 259018 509946 259254
rect 510182 259018 510266 259254
rect 510502 259018 510534 259254
rect 509914 223574 510534 259018
rect 509914 223338 509946 223574
rect 510182 223338 510266 223574
rect 510502 223338 510534 223574
rect 509914 223254 510534 223338
rect 509914 223018 509946 223254
rect 510182 223018 510266 223254
rect 510502 223018 510534 223254
rect 509914 187574 510534 223018
rect 509914 187338 509946 187574
rect 510182 187338 510266 187574
rect 510502 187338 510534 187574
rect 509914 187254 510534 187338
rect 509914 187018 509946 187254
rect 510182 187018 510266 187254
rect 510502 187018 510534 187254
rect 509914 151574 510534 187018
rect 509914 151338 509946 151574
rect 510182 151338 510266 151574
rect 510502 151338 510534 151574
rect 509914 151254 510534 151338
rect 509914 151018 509946 151254
rect 510182 151018 510266 151254
rect 510502 151018 510534 151254
rect 509914 115574 510534 151018
rect 509914 115338 509946 115574
rect 510182 115338 510266 115574
rect 510502 115338 510534 115574
rect 509914 115254 510534 115338
rect 509914 115018 509946 115254
rect 510182 115018 510266 115254
rect 510502 115018 510534 115254
rect 509914 79574 510534 115018
rect 509914 79338 509946 79574
rect 510182 79338 510266 79574
rect 510502 79338 510534 79574
rect 509914 79254 510534 79338
rect 509914 79018 509946 79254
rect 510182 79018 510266 79254
rect 510502 79018 510534 79254
rect 509914 43574 510534 79018
rect 509914 43338 509946 43574
rect 510182 43338 510266 43574
rect 510502 43338 510534 43574
rect 509914 43254 510534 43338
rect 509914 43018 509946 43254
rect 510182 43018 510266 43254
rect 510502 43018 510534 43254
rect 509914 7574 510534 43018
rect 509914 7338 509946 7574
rect 510182 7338 510266 7574
rect 510502 7338 510534 7574
rect 509914 7254 510534 7338
rect 509914 7018 509946 7254
rect 510182 7018 510266 7254
rect 510502 7018 510534 7254
rect 509914 -1306 510534 7018
rect 509914 -1542 509946 -1306
rect 510182 -1542 510266 -1306
rect 510502 -1542 510534 -1306
rect 509914 -1626 510534 -1542
rect 509914 -1862 509946 -1626
rect 510182 -1862 510266 -1626
rect 510502 -1862 510534 -1626
rect 509914 -7654 510534 -1862
rect 513634 706758 514254 711590
rect 513634 706522 513666 706758
rect 513902 706522 513986 706758
rect 514222 706522 514254 706758
rect 513634 706438 514254 706522
rect 513634 706202 513666 706438
rect 513902 706202 513986 706438
rect 514222 706202 514254 706438
rect 513634 695294 514254 706202
rect 513634 695058 513666 695294
rect 513902 695058 513986 695294
rect 514222 695058 514254 695294
rect 513634 694974 514254 695058
rect 513634 694738 513666 694974
rect 513902 694738 513986 694974
rect 514222 694738 514254 694974
rect 513634 659294 514254 694738
rect 513634 659058 513666 659294
rect 513902 659058 513986 659294
rect 514222 659058 514254 659294
rect 513634 658974 514254 659058
rect 513634 658738 513666 658974
rect 513902 658738 513986 658974
rect 514222 658738 514254 658974
rect 513634 623294 514254 658738
rect 513634 623058 513666 623294
rect 513902 623058 513986 623294
rect 514222 623058 514254 623294
rect 513634 622974 514254 623058
rect 513634 622738 513666 622974
rect 513902 622738 513986 622974
rect 514222 622738 514254 622974
rect 513634 587294 514254 622738
rect 513634 587058 513666 587294
rect 513902 587058 513986 587294
rect 514222 587058 514254 587294
rect 513634 586974 514254 587058
rect 513634 586738 513666 586974
rect 513902 586738 513986 586974
rect 514222 586738 514254 586974
rect 513634 551294 514254 586738
rect 513634 551058 513666 551294
rect 513902 551058 513986 551294
rect 514222 551058 514254 551294
rect 513634 550974 514254 551058
rect 513634 550738 513666 550974
rect 513902 550738 513986 550974
rect 514222 550738 514254 550974
rect 513634 515294 514254 550738
rect 513634 515058 513666 515294
rect 513902 515058 513986 515294
rect 514222 515058 514254 515294
rect 513634 514974 514254 515058
rect 513634 514738 513666 514974
rect 513902 514738 513986 514974
rect 514222 514738 514254 514974
rect 513634 479294 514254 514738
rect 513634 479058 513666 479294
rect 513902 479058 513986 479294
rect 514222 479058 514254 479294
rect 513634 478974 514254 479058
rect 513634 478738 513666 478974
rect 513902 478738 513986 478974
rect 514222 478738 514254 478974
rect 513634 443294 514254 478738
rect 513634 443058 513666 443294
rect 513902 443058 513986 443294
rect 514222 443058 514254 443294
rect 513634 442974 514254 443058
rect 513634 442738 513666 442974
rect 513902 442738 513986 442974
rect 514222 442738 514254 442974
rect 513634 407294 514254 442738
rect 513634 407058 513666 407294
rect 513902 407058 513986 407294
rect 514222 407058 514254 407294
rect 513634 406974 514254 407058
rect 513634 406738 513666 406974
rect 513902 406738 513986 406974
rect 514222 406738 514254 406974
rect 513634 371294 514254 406738
rect 513634 371058 513666 371294
rect 513902 371058 513986 371294
rect 514222 371058 514254 371294
rect 513634 370974 514254 371058
rect 513634 370738 513666 370974
rect 513902 370738 513986 370974
rect 514222 370738 514254 370974
rect 513634 335294 514254 370738
rect 513634 335058 513666 335294
rect 513902 335058 513986 335294
rect 514222 335058 514254 335294
rect 513634 334974 514254 335058
rect 513634 334738 513666 334974
rect 513902 334738 513986 334974
rect 514222 334738 514254 334974
rect 513634 299294 514254 334738
rect 513634 299058 513666 299294
rect 513902 299058 513986 299294
rect 514222 299058 514254 299294
rect 513634 298974 514254 299058
rect 513634 298738 513666 298974
rect 513902 298738 513986 298974
rect 514222 298738 514254 298974
rect 513634 263294 514254 298738
rect 513634 263058 513666 263294
rect 513902 263058 513986 263294
rect 514222 263058 514254 263294
rect 513634 262974 514254 263058
rect 513634 262738 513666 262974
rect 513902 262738 513986 262974
rect 514222 262738 514254 262974
rect 513634 227294 514254 262738
rect 513634 227058 513666 227294
rect 513902 227058 513986 227294
rect 514222 227058 514254 227294
rect 513634 226974 514254 227058
rect 513634 226738 513666 226974
rect 513902 226738 513986 226974
rect 514222 226738 514254 226974
rect 513634 191294 514254 226738
rect 513634 191058 513666 191294
rect 513902 191058 513986 191294
rect 514222 191058 514254 191294
rect 513634 190974 514254 191058
rect 513634 190738 513666 190974
rect 513902 190738 513986 190974
rect 514222 190738 514254 190974
rect 513634 155294 514254 190738
rect 513634 155058 513666 155294
rect 513902 155058 513986 155294
rect 514222 155058 514254 155294
rect 513634 154974 514254 155058
rect 513634 154738 513666 154974
rect 513902 154738 513986 154974
rect 514222 154738 514254 154974
rect 513634 119294 514254 154738
rect 513634 119058 513666 119294
rect 513902 119058 513986 119294
rect 514222 119058 514254 119294
rect 513634 118974 514254 119058
rect 513634 118738 513666 118974
rect 513902 118738 513986 118974
rect 514222 118738 514254 118974
rect 513634 83294 514254 118738
rect 513634 83058 513666 83294
rect 513902 83058 513986 83294
rect 514222 83058 514254 83294
rect 513634 82974 514254 83058
rect 513634 82738 513666 82974
rect 513902 82738 513986 82974
rect 514222 82738 514254 82974
rect 513634 47294 514254 82738
rect 513634 47058 513666 47294
rect 513902 47058 513986 47294
rect 514222 47058 514254 47294
rect 513634 46974 514254 47058
rect 513634 46738 513666 46974
rect 513902 46738 513986 46974
rect 514222 46738 514254 46974
rect 513634 11294 514254 46738
rect 513634 11058 513666 11294
rect 513902 11058 513986 11294
rect 514222 11058 514254 11294
rect 513634 10974 514254 11058
rect 513634 10738 513666 10974
rect 513902 10738 513986 10974
rect 514222 10738 514254 10974
rect 513634 -2266 514254 10738
rect 513634 -2502 513666 -2266
rect 513902 -2502 513986 -2266
rect 514222 -2502 514254 -2266
rect 513634 -2586 514254 -2502
rect 513634 -2822 513666 -2586
rect 513902 -2822 513986 -2586
rect 514222 -2822 514254 -2586
rect 513634 -7654 514254 -2822
rect 517354 707718 517974 711590
rect 517354 707482 517386 707718
rect 517622 707482 517706 707718
rect 517942 707482 517974 707718
rect 517354 707398 517974 707482
rect 517354 707162 517386 707398
rect 517622 707162 517706 707398
rect 517942 707162 517974 707398
rect 517354 699014 517974 707162
rect 517354 698778 517386 699014
rect 517622 698778 517706 699014
rect 517942 698778 517974 699014
rect 517354 698694 517974 698778
rect 517354 698458 517386 698694
rect 517622 698458 517706 698694
rect 517942 698458 517974 698694
rect 517354 663014 517974 698458
rect 517354 662778 517386 663014
rect 517622 662778 517706 663014
rect 517942 662778 517974 663014
rect 517354 662694 517974 662778
rect 517354 662458 517386 662694
rect 517622 662458 517706 662694
rect 517942 662458 517974 662694
rect 517354 627014 517974 662458
rect 517354 626778 517386 627014
rect 517622 626778 517706 627014
rect 517942 626778 517974 627014
rect 517354 626694 517974 626778
rect 517354 626458 517386 626694
rect 517622 626458 517706 626694
rect 517942 626458 517974 626694
rect 517354 591014 517974 626458
rect 517354 590778 517386 591014
rect 517622 590778 517706 591014
rect 517942 590778 517974 591014
rect 517354 590694 517974 590778
rect 517354 590458 517386 590694
rect 517622 590458 517706 590694
rect 517942 590458 517974 590694
rect 517354 555014 517974 590458
rect 517354 554778 517386 555014
rect 517622 554778 517706 555014
rect 517942 554778 517974 555014
rect 517354 554694 517974 554778
rect 517354 554458 517386 554694
rect 517622 554458 517706 554694
rect 517942 554458 517974 554694
rect 517354 519014 517974 554458
rect 517354 518778 517386 519014
rect 517622 518778 517706 519014
rect 517942 518778 517974 519014
rect 517354 518694 517974 518778
rect 517354 518458 517386 518694
rect 517622 518458 517706 518694
rect 517942 518458 517974 518694
rect 517354 483014 517974 518458
rect 517354 482778 517386 483014
rect 517622 482778 517706 483014
rect 517942 482778 517974 483014
rect 517354 482694 517974 482778
rect 517354 482458 517386 482694
rect 517622 482458 517706 482694
rect 517942 482458 517974 482694
rect 517354 447014 517974 482458
rect 517354 446778 517386 447014
rect 517622 446778 517706 447014
rect 517942 446778 517974 447014
rect 517354 446694 517974 446778
rect 517354 446458 517386 446694
rect 517622 446458 517706 446694
rect 517942 446458 517974 446694
rect 517354 411014 517974 446458
rect 517354 410778 517386 411014
rect 517622 410778 517706 411014
rect 517942 410778 517974 411014
rect 517354 410694 517974 410778
rect 517354 410458 517386 410694
rect 517622 410458 517706 410694
rect 517942 410458 517974 410694
rect 517354 375014 517974 410458
rect 517354 374778 517386 375014
rect 517622 374778 517706 375014
rect 517942 374778 517974 375014
rect 517354 374694 517974 374778
rect 517354 374458 517386 374694
rect 517622 374458 517706 374694
rect 517942 374458 517974 374694
rect 517354 339014 517974 374458
rect 517354 338778 517386 339014
rect 517622 338778 517706 339014
rect 517942 338778 517974 339014
rect 517354 338694 517974 338778
rect 517354 338458 517386 338694
rect 517622 338458 517706 338694
rect 517942 338458 517974 338694
rect 517354 303014 517974 338458
rect 517354 302778 517386 303014
rect 517622 302778 517706 303014
rect 517942 302778 517974 303014
rect 517354 302694 517974 302778
rect 517354 302458 517386 302694
rect 517622 302458 517706 302694
rect 517942 302458 517974 302694
rect 517354 267014 517974 302458
rect 517354 266778 517386 267014
rect 517622 266778 517706 267014
rect 517942 266778 517974 267014
rect 517354 266694 517974 266778
rect 517354 266458 517386 266694
rect 517622 266458 517706 266694
rect 517942 266458 517974 266694
rect 517354 231014 517974 266458
rect 517354 230778 517386 231014
rect 517622 230778 517706 231014
rect 517942 230778 517974 231014
rect 517354 230694 517974 230778
rect 517354 230458 517386 230694
rect 517622 230458 517706 230694
rect 517942 230458 517974 230694
rect 517354 195014 517974 230458
rect 517354 194778 517386 195014
rect 517622 194778 517706 195014
rect 517942 194778 517974 195014
rect 517354 194694 517974 194778
rect 517354 194458 517386 194694
rect 517622 194458 517706 194694
rect 517942 194458 517974 194694
rect 517354 159014 517974 194458
rect 517354 158778 517386 159014
rect 517622 158778 517706 159014
rect 517942 158778 517974 159014
rect 517354 158694 517974 158778
rect 517354 158458 517386 158694
rect 517622 158458 517706 158694
rect 517942 158458 517974 158694
rect 517354 123014 517974 158458
rect 517354 122778 517386 123014
rect 517622 122778 517706 123014
rect 517942 122778 517974 123014
rect 517354 122694 517974 122778
rect 517354 122458 517386 122694
rect 517622 122458 517706 122694
rect 517942 122458 517974 122694
rect 517354 87014 517974 122458
rect 517354 86778 517386 87014
rect 517622 86778 517706 87014
rect 517942 86778 517974 87014
rect 517354 86694 517974 86778
rect 517354 86458 517386 86694
rect 517622 86458 517706 86694
rect 517942 86458 517974 86694
rect 517354 51014 517974 86458
rect 517354 50778 517386 51014
rect 517622 50778 517706 51014
rect 517942 50778 517974 51014
rect 517354 50694 517974 50778
rect 517354 50458 517386 50694
rect 517622 50458 517706 50694
rect 517942 50458 517974 50694
rect 517354 15014 517974 50458
rect 517354 14778 517386 15014
rect 517622 14778 517706 15014
rect 517942 14778 517974 15014
rect 517354 14694 517974 14778
rect 517354 14458 517386 14694
rect 517622 14458 517706 14694
rect 517942 14458 517974 14694
rect 517354 -3226 517974 14458
rect 517354 -3462 517386 -3226
rect 517622 -3462 517706 -3226
rect 517942 -3462 517974 -3226
rect 517354 -3546 517974 -3462
rect 517354 -3782 517386 -3546
rect 517622 -3782 517706 -3546
rect 517942 -3782 517974 -3546
rect 517354 -7654 517974 -3782
rect 521074 708678 521694 711590
rect 521074 708442 521106 708678
rect 521342 708442 521426 708678
rect 521662 708442 521694 708678
rect 521074 708358 521694 708442
rect 521074 708122 521106 708358
rect 521342 708122 521426 708358
rect 521662 708122 521694 708358
rect 521074 666734 521694 708122
rect 521074 666498 521106 666734
rect 521342 666498 521426 666734
rect 521662 666498 521694 666734
rect 521074 666414 521694 666498
rect 521074 666178 521106 666414
rect 521342 666178 521426 666414
rect 521662 666178 521694 666414
rect 521074 630734 521694 666178
rect 521074 630498 521106 630734
rect 521342 630498 521426 630734
rect 521662 630498 521694 630734
rect 521074 630414 521694 630498
rect 521074 630178 521106 630414
rect 521342 630178 521426 630414
rect 521662 630178 521694 630414
rect 521074 594734 521694 630178
rect 521074 594498 521106 594734
rect 521342 594498 521426 594734
rect 521662 594498 521694 594734
rect 521074 594414 521694 594498
rect 521074 594178 521106 594414
rect 521342 594178 521426 594414
rect 521662 594178 521694 594414
rect 521074 558734 521694 594178
rect 521074 558498 521106 558734
rect 521342 558498 521426 558734
rect 521662 558498 521694 558734
rect 521074 558414 521694 558498
rect 521074 558178 521106 558414
rect 521342 558178 521426 558414
rect 521662 558178 521694 558414
rect 521074 522734 521694 558178
rect 521074 522498 521106 522734
rect 521342 522498 521426 522734
rect 521662 522498 521694 522734
rect 521074 522414 521694 522498
rect 521074 522178 521106 522414
rect 521342 522178 521426 522414
rect 521662 522178 521694 522414
rect 521074 486734 521694 522178
rect 521074 486498 521106 486734
rect 521342 486498 521426 486734
rect 521662 486498 521694 486734
rect 521074 486414 521694 486498
rect 521074 486178 521106 486414
rect 521342 486178 521426 486414
rect 521662 486178 521694 486414
rect 521074 450734 521694 486178
rect 521074 450498 521106 450734
rect 521342 450498 521426 450734
rect 521662 450498 521694 450734
rect 521074 450414 521694 450498
rect 521074 450178 521106 450414
rect 521342 450178 521426 450414
rect 521662 450178 521694 450414
rect 521074 414734 521694 450178
rect 521074 414498 521106 414734
rect 521342 414498 521426 414734
rect 521662 414498 521694 414734
rect 521074 414414 521694 414498
rect 521074 414178 521106 414414
rect 521342 414178 521426 414414
rect 521662 414178 521694 414414
rect 521074 378734 521694 414178
rect 521074 378498 521106 378734
rect 521342 378498 521426 378734
rect 521662 378498 521694 378734
rect 521074 378414 521694 378498
rect 521074 378178 521106 378414
rect 521342 378178 521426 378414
rect 521662 378178 521694 378414
rect 521074 342734 521694 378178
rect 521074 342498 521106 342734
rect 521342 342498 521426 342734
rect 521662 342498 521694 342734
rect 521074 342414 521694 342498
rect 521074 342178 521106 342414
rect 521342 342178 521426 342414
rect 521662 342178 521694 342414
rect 521074 306734 521694 342178
rect 521074 306498 521106 306734
rect 521342 306498 521426 306734
rect 521662 306498 521694 306734
rect 521074 306414 521694 306498
rect 521074 306178 521106 306414
rect 521342 306178 521426 306414
rect 521662 306178 521694 306414
rect 521074 270734 521694 306178
rect 521074 270498 521106 270734
rect 521342 270498 521426 270734
rect 521662 270498 521694 270734
rect 521074 270414 521694 270498
rect 521074 270178 521106 270414
rect 521342 270178 521426 270414
rect 521662 270178 521694 270414
rect 521074 234734 521694 270178
rect 521074 234498 521106 234734
rect 521342 234498 521426 234734
rect 521662 234498 521694 234734
rect 521074 234414 521694 234498
rect 521074 234178 521106 234414
rect 521342 234178 521426 234414
rect 521662 234178 521694 234414
rect 521074 198734 521694 234178
rect 521074 198498 521106 198734
rect 521342 198498 521426 198734
rect 521662 198498 521694 198734
rect 521074 198414 521694 198498
rect 521074 198178 521106 198414
rect 521342 198178 521426 198414
rect 521662 198178 521694 198414
rect 521074 162734 521694 198178
rect 521074 162498 521106 162734
rect 521342 162498 521426 162734
rect 521662 162498 521694 162734
rect 521074 162414 521694 162498
rect 521074 162178 521106 162414
rect 521342 162178 521426 162414
rect 521662 162178 521694 162414
rect 521074 126734 521694 162178
rect 521074 126498 521106 126734
rect 521342 126498 521426 126734
rect 521662 126498 521694 126734
rect 521074 126414 521694 126498
rect 521074 126178 521106 126414
rect 521342 126178 521426 126414
rect 521662 126178 521694 126414
rect 521074 90734 521694 126178
rect 521074 90498 521106 90734
rect 521342 90498 521426 90734
rect 521662 90498 521694 90734
rect 521074 90414 521694 90498
rect 521074 90178 521106 90414
rect 521342 90178 521426 90414
rect 521662 90178 521694 90414
rect 521074 54734 521694 90178
rect 521074 54498 521106 54734
rect 521342 54498 521426 54734
rect 521662 54498 521694 54734
rect 521074 54414 521694 54498
rect 521074 54178 521106 54414
rect 521342 54178 521426 54414
rect 521662 54178 521694 54414
rect 521074 18734 521694 54178
rect 521074 18498 521106 18734
rect 521342 18498 521426 18734
rect 521662 18498 521694 18734
rect 521074 18414 521694 18498
rect 521074 18178 521106 18414
rect 521342 18178 521426 18414
rect 521662 18178 521694 18414
rect 521074 -4186 521694 18178
rect 521074 -4422 521106 -4186
rect 521342 -4422 521426 -4186
rect 521662 -4422 521694 -4186
rect 521074 -4506 521694 -4422
rect 521074 -4742 521106 -4506
rect 521342 -4742 521426 -4506
rect 521662 -4742 521694 -4506
rect 521074 -7654 521694 -4742
rect 524794 709638 525414 711590
rect 524794 709402 524826 709638
rect 525062 709402 525146 709638
rect 525382 709402 525414 709638
rect 524794 709318 525414 709402
rect 524794 709082 524826 709318
rect 525062 709082 525146 709318
rect 525382 709082 525414 709318
rect 524794 670454 525414 709082
rect 524794 670218 524826 670454
rect 525062 670218 525146 670454
rect 525382 670218 525414 670454
rect 524794 670134 525414 670218
rect 524794 669898 524826 670134
rect 525062 669898 525146 670134
rect 525382 669898 525414 670134
rect 524794 634454 525414 669898
rect 524794 634218 524826 634454
rect 525062 634218 525146 634454
rect 525382 634218 525414 634454
rect 524794 634134 525414 634218
rect 524794 633898 524826 634134
rect 525062 633898 525146 634134
rect 525382 633898 525414 634134
rect 524794 598454 525414 633898
rect 524794 598218 524826 598454
rect 525062 598218 525146 598454
rect 525382 598218 525414 598454
rect 524794 598134 525414 598218
rect 524794 597898 524826 598134
rect 525062 597898 525146 598134
rect 525382 597898 525414 598134
rect 524794 562454 525414 597898
rect 524794 562218 524826 562454
rect 525062 562218 525146 562454
rect 525382 562218 525414 562454
rect 524794 562134 525414 562218
rect 524794 561898 524826 562134
rect 525062 561898 525146 562134
rect 525382 561898 525414 562134
rect 524794 526454 525414 561898
rect 524794 526218 524826 526454
rect 525062 526218 525146 526454
rect 525382 526218 525414 526454
rect 524794 526134 525414 526218
rect 524794 525898 524826 526134
rect 525062 525898 525146 526134
rect 525382 525898 525414 526134
rect 524794 490454 525414 525898
rect 524794 490218 524826 490454
rect 525062 490218 525146 490454
rect 525382 490218 525414 490454
rect 524794 490134 525414 490218
rect 524794 489898 524826 490134
rect 525062 489898 525146 490134
rect 525382 489898 525414 490134
rect 524794 454454 525414 489898
rect 524794 454218 524826 454454
rect 525062 454218 525146 454454
rect 525382 454218 525414 454454
rect 524794 454134 525414 454218
rect 524794 453898 524826 454134
rect 525062 453898 525146 454134
rect 525382 453898 525414 454134
rect 524794 418454 525414 453898
rect 524794 418218 524826 418454
rect 525062 418218 525146 418454
rect 525382 418218 525414 418454
rect 524794 418134 525414 418218
rect 524794 417898 524826 418134
rect 525062 417898 525146 418134
rect 525382 417898 525414 418134
rect 524794 382454 525414 417898
rect 524794 382218 524826 382454
rect 525062 382218 525146 382454
rect 525382 382218 525414 382454
rect 524794 382134 525414 382218
rect 524794 381898 524826 382134
rect 525062 381898 525146 382134
rect 525382 381898 525414 382134
rect 524794 346454 525414 381898
rect 524794 346218 524826 346454
rect 525062 346218 525146 346454
rect 525382 346218 525414 346454
rect 524794 346134 525414 346218
rect 524794 345898 524826 346134
rect 525062 345898 525146 346134
rect 525382 345898 525414 346134
rect 524794 310454 525414 345898
rect 524794 310218 524826 310454
rect 525062 310218 525146 310454
rect 525382 310218 525414 310454
rect 524794 310134 525414 310218
rect 524794 309898 524826 310134
rect 525062 309898 525146 310134
rect 525382 309898 525414 310134
rect 524794 274454 525414 309898
rect 524794 274218 524826 274454
rect 525062 274218 525146 274454
rect 525382 274218 525414 274454
rect 524794 274134 525414 274218
rect 524794 273898 524826 274134
rect 525062 273898 525146 274134
rect 525382 273898 525414 274134
rect 524794 238454 525414 273898
rect 524794 238218 524826 238454
rect 525062 238218 525146 238454
rect 525382 238218 525414 238454
rect 524794 238134 525414 238218
rect 524794 237898 524826 238134
rect 525062 237898 525146 238134
rect 525382 237898 525414 238134
rect 524794 202454 525414 237898
rect 524794 202218 524826 202454
rect 525062 202218 525146 202454
rect 525382 202218 525414 202454
rect 524794 202134 525414 202218
rect 524794 201898 524826 202134
rect 525062 201898 525146 202134
rect 525382 201898 525414 202134
rect 524794 166454 525414 201898
rect 524794 166218 524826 166454
rect 525062 166218 525146 166454
rect 525382 166218 525414 166454
rect 524794 166134 525414 166218
rect 524794 165898 524826 166134
rect 525062 165898 525146 166134
rect 525382 165898 525414 166134
rect 524794 130454 525414 165898
rect 524794 130218 524826 130454
rect 525062 130218 525146 130454
rect 525382 130218 525414 130454
rect 524794 130134 525414 130218
rect 524794 129898 524826 130134
rect 525062 129898 525146 130134
rect 525382 129898 525414 130134
rect 524794 94454 525414 129898
rect 524794 94218 524826 94454
rect 525062 94218 525146 94454
rect 525382 94218 525414 94454
rect 524794 94134 525414 94218
rect 524794 93898 524826 94134
rect 525062 93898 525146 94134
rect 525382 93898 525414 94134
rect 524794 58454 525414 93898
rect 524794 58218 524826 58454
rect 525062 58218 525146 58454
rect 525382 58218 525414 58454
rect 524794 58134 525414 58218
rect 524794 57898 524826 58134
rect 525062 57898 525146 58134
rect 525382 57898 525414 58134
rect 524794 22454 525414 57898
rect 524794 22218 524826 22454
rect 525062 22218 525146 22454
rect 525382 22218 525414 22454
rect 524794 22134 525414 22218
rect 524794 21898 524826 22134
rect 525062 21898 525146 22134
rect 525382 21898 525414 22134
rect 524794 -5146 525414 21898
rect 524794 -5382 524826 -5146
rect 525062 -5382 525146 -5146
rect 525382 -5382 525414 -5146
rect 524794 -5466 525414 -5382
rect 524794 -5702 524826 -5466
rect 525062 -5702 525146 -5466
rect 525382 -5702 525414 -5466
rect 524794 -7654 525414 -5702
rect 528514 710598 529134 711590
rect 528514 710362 528546 710598
rect 528782 710362 528866 710598
rect 529102 710362 529134 710598
rect 528514 710278 529134 710362
rect 528514 710042 528546 710278
rect 528782 710042 528866 710278
rect 529102 710042 529134 710278
rect 528514 674174 529134 710042
rect 528514 673938 528546 674174
rect 528782 673938 528866 674174
rect 529102 673938 529134 674174
rect 528514 673854 529134 673938
rect 528514 673618 528546 673854
rect 528782 673618 528866 673854
rect 529102 673618 529134 673854
rect 528514 638174 529134 673618
rect 528514 637938 528546 638174
rect 528782 637938 528866 638174
rect 529102 637938 529134 638174
rect 528514 637854 529134 637938
rect 528514 637618 528546 637854
rect 528782 637618 528866 637854
rect 529102 637618 529134 637854
rect 528514 602174 529134 637618
rect 528514 601938 528546 602174
rect 528782 601938 528866 602174
rect 529102 601938 529134 602174
rect 528514 601854 529134 601938
rect 528514 601618 528546 601854
rect 528782 601618 528866 601854
rect 529102 601618 529134 601854
rect 528514 566174 529134 601618
rect 528514 565938 528546 566174
rect 528782 565938 528866 566174
rect 529102 565938 529134 566174
rect 528514 565854 529134 565938
rect 528514 565618 528546 565854
rect 528782 565618 528866 565854
rect 529102 565618 529134 565854
rect 528514 530174 529134 565618
rect 528514 529938 528546 530174
rect 528782 529938 528866 530174
rect 529102 529938 529134 530174
rect 528514 529854 529134 529938
rect 528514 529618 528546 529854
rect 528782 529618 528866 529854
rect 529102 529618 529134 529854
rect 528514 494174 529134 529618
rect 528514 493938 528546 494174
rect 528782 493938 528866 494174
rect 529102 493938 529134 494174
rect 528514 493854 529134 493938
rect 528514 493618 528546 493854
rect 528782 493618 528866 493854
rect 529102 493618 529134 493854
rect 528514 458174 529134 493618
rect 528514 457938 528546 458174
rect 528782 457938 528866 458174
rect 529102 457938 529134 458174
rect 528514 457854 529134 457938
rect 528514 457618 528546 457854
rect 528782 457618 528866 457854
rect 529102 457618 529134 457854
rect 528514 422174 529134 457618
rect 528514 421938 528546 422174
rect 528782 421938 528866 422174
rect 529102 421938 529134 422174
rect 528514 421854 529134 421938
rect 528514 421618 528546 421854
rect 528782 421618 528866 421854
rect 529102 421618 529134 421854
rect 528514 386174 529134 421618
rect 528514 385938 528546 386174
rect 528782 385938 528866 386174
rect 529102 385938 529134 386174
rect 528514 385854 529134 385938
rect 528514 385618 528546 385854
rect 528782 385618 528866 385854
rect 529102 385618 529134 385854
rect 528514 350174 529134 385618
rect 528514 349938 528546 350174
rect 528782 349938 528866 350174
rect 529102 349938 529134 350174
rect 528514 349854 529134 349938
rect 528514 349618 528546 349854
rect 528782 349618 528866 349854
rect 529102 349618 529134 349854
rect 528514 314174 529134 349618
rect 528514 313938 528546 314174
rect 528782 313938 528866 314174
rect 529102 313938 529134 314174
rect 528514 313854 529134 313938
rect 528514 313618 528546 313854
rect 528782 313618 528866 313854
rect 529102 313618 529134 313854
rect 528514 278174 529134 313618
rect 528514 277938 528546 278174
rect 528782 277938 528866 278174
rect 529102 277938 529134 278174
rect 528514 277854 529134 277938
rect 528514 277618 528546 277854
rect 528782 277618 528866 277854
rect 529102 277618 529134 277854
rect 528514 242174 529134 277618
rect 528514 241938 528546 242174
rect 528782 241938 528866 242174
rect 529102 241938 529134 242174
rect 528514 241854 529134 241938
rect 528514 241618 528546 241854
rect 528782 241618 528866 241854
rect 529102 241618 529134 241854
rect 528514 206174 529134 241618
rect 528514 205938 528546 206174
rect 528782 205938 528866 206174
rect 529102 205938 529134 206174
rect 528514 205854 529134 205938
rect 528514 205618 528546 205854
rect 528782 205618 528866 205854
rect 529102 205618 529134 205854
rect 528514 170174 529134 205618
rect 528514 169938 528546 170174
rect 528782 169938 528866 170174
rect 529102 169938 529134 170174
rect 528514 169854 529134 169938
rect 528514 169618 528546 169854
rect 528782 169618 528866 169854
rect 529102 169618 529134 169854
rect 528514 134174 529134 169618
rect 528514 133938 528546 134174
rect 528782 133938 528866 134174
rect 529102 133938 529134 134174
rect 528514 133854 529134 133938
rect 528514 133618 528546 133854
rect 528782 133618 528866 133854
rect 529102 133618 529134 133854
rect 528514 98174 529134 133618
rect 528514 97938 528546 98174
rect 528782 97938 528866 98174
rect 529102 97938 529134 98174
rect 528514 97854 529134 97938
rect 528514 97618 528546 97854
rect 528782 97618 528866 97854
rect 529102 97618 529134 97854
rect 528514 62174 529134 97618
rect 528514 61938 528546 62174
rect 528782 61938 528866 62174
rect 529102 61938 529134 62174
rect 528514 61854 529134 61938
rect 528514 61618 528546 61854
rect 528782 61618 528866 61854
rect 529102 61618 529134 61854
rect 528514 26174 529134 61618
rect 528514 25938 528546 26174
rect 528782 25938 528866 26174
rect 529102 25938 529134 26174
rect 528514 25854 529134 25938
rect 528514 25618 528546 25854
rect 528782 25618 528866 25854
rect 529102 25618 529134 25854
rect 528514 -6106 529134 25618
rect 528514 -6342 528546 -6106
rect 528782 -6342 528866 -6106
rect 529102 -6342 529134 -6106
rect 528514 -6426 529134 -6342
rect 528514 -6662 528546 -6426
rect 528782 -6662 528866 -6426
rect 529102 -6662 529134 -6426
rect 528514 -7654 529134 -6662
rect 532234 711558 532854 711590
rect 532234 711322 532266 711558
rect 532502 711322 532586 711558
rect 532822 711322 532854 711558
rect 532234 711238 532854 711322
rect 532234 711002 532266 711238
rect 532502 711002 532586 711238
rect 532822 711002 532854 711238
rect 532234 677894 532854 711002
rect 532234 677658 532266 677894
rect 532502 677658 532586 677894
rect 532822 677658 532854 677894
rect 532234 677574 532854 677658
rect 532234 677338 532266 677574
rect 532502 677338 532586 677574
rect 532822 677338 532854 677574
rect 532234 641894 532854 677338
rect 532234 641658 532266 641894
rect 532502 641658 532586 641894
rect 532822 641658 532854 641894
rect 532234 641574 532854 641658
rect 532234 641338 532266 641574
rect 532502 641338 532586 641574
rect 532822 641338 532854 641574
rect 532234 605894 532854 641338
rect 532234 605658 532266 605894
rect 532502 605658 532586 605894
rect 532822 605658 532854 605894
rect 532234 605574 532854 605658
rect 532234 605338 532266 605574
rect 532502 605338 532586 605574
rect 532822 605338 532854 605574
rect 532234 569894 532854 605338
rect 532234 569658 532266 569894
rect 532502 569658 532586 569894
rect 532822 569658 532854 569894
rect 532234 569574 532854 569658
rect 532234 569338 532266 569574
rect 532502 569338 532586 569574
rect 532822 569338 532854 569574
rect 532234 533894 532854 569338
rect 532234 533658 532266 533894
rect 532502 533658 532586 533894
rect 532822 533658 532854 533894
rect 532234 533574 532854 533658
rect 532234 533338 532266 533574
rect 532502 533338 532586 533574
rect 532822 533338 532854 533574
rect 532234 497894 532854 533338
rect 532234 497658 532266 497894
rect 532502 497658 532586 497894
rect 532822 497658 532854 497894
rect 532234 497574 532854 497658
rect 532234 497338 532266 497574
rect 532502 497338 532586 497574
rect 532822 497338 532854 497574
rect 532234 461894 532854 497338
rect 532234 461658 532266 461894
rect 532502 461658 532586 461894
rect 532822 461658 532854 461894
rect 532234 461574 532854 461658
rect 532234 461338 532266 461574
rect 532502 461338 532586 461574
rect 532822 461338 532854 461574
rect 532234 425894 532854 461338
rect 532234 425658 532266 425894
rect 532502 425658 532586 425894
rect 532822 425658 532854 425894
rect 532234 425574 532854 425658
rect 532234 425338 532266 425574
rect 532502 425338 532586 425574
rect 532822 425338 532854 425574
rect 532234 389894 532854 425338
rect 532234 389658 532266 389894
rect 532502 389658 532586 389894
rect 532822 389658 532854 389894
rect 532234 389574 532854 389658
rect 532234 389338 532266 389574
rect 532502 389338 532586 389574
rect 532822 389338 532854 389574
rect 532234 353894 532854 389338
rect 532234 353658 532266 353894
rect 532502 353658 532586 353894
rect 532822 353658 532854 353894
rect 532234 353574 532854 353658
rect 532234 353338 532266 353574
rect 532502 353338 532586 353574
rect 532822 353338 532854 353574
rect 532234 317894 532854 353338
rect 532234 317658 532266 317894
rect 532502 317658 532586 317894
rect 532822 317658 532854 317894
rect 532234 317574 532854 317658
rect 532234 317338 532266 317574
rect 532502 317338 532586 317574
rect 532822 317338 532854 317574
rect 532234 281894 532854 317338
rect 532234 281658 532266 281894
rect 532502 281658 532586 281894
rect 532822 281658 532854 281894
rect 532234 281574 532854 281658
rect 532234 281338 532266 281574
rect 532502 281338 532586 281574
rect 532822 281338 532854 281574
rect 532234 245894 532854 281338
rect 532234 245658 532266 245894
rect 532502 245658 532586 245894
rect 532822 245658 532854 245894
rect 532234 245574 532854 245658
rect 532234 245338 532266 245574
rect 532502 245338 532586 245574
rect 532822 245338 532854 245574
rect 532234 209894 532854 245338
rect 532234 209658 532266 209894
rect 532502 209658 532586 209894
rect 532822 209658 532854 209894
rect 532234 209574 532854 209658
rect 532234 209338 532266 209574
rect 532502 209338 532586 209574
rect 532822 209338 532854 209574
rect 532234 173894 532854 209338
rect 532234 173658 532266 173894
rect 532502 173658 532586 173894
rect 532822 173658 532854 173894
rect 532234 173574 532854 173658
rect 532234 173338 532266 173574
rect 532502 173338 532586 173574
rect 532822 173338 532854 173574
rect 532234 137894 532854 173338
rect 532234 137658 532266 137894
rect 532502 137658 532586 137894
rect 532822 137658 532854 137894
rect 532234 137574 532854 137658
rect 532234 137338 532266 137574
rect 532502 137338 532586 137574
rect 532822 137338 532854 137574
rect 532234 101894 532854 137338
rect 532234 101658 532266 101894
rect 532502 101658 532586 101894
rect 532822 101658 532854 101894
rect 532234 101574 532854 101658
rect 532234 101338 532266 101574
rect 532502 101338 532586 101574
rect 532822 101338 532854 101574
rect 532234 65894 532854 101338
rect 532234 65658 532266 65894
rect 532502 65658 532586 65894
rect 532822 65658 532854 65894
rect 532234 65574 532854 65658
rect 532234 65338 532266 65574
rect 532502 65338 532586 65574
rect 532822 65338 532854 65574
rect 532234 29894 532854 65338
rect 532234 29658 532266 29894
rect 532502 29658 532586 29894
rect 532822 29658 532854 29894
rect 532234 29574 532854 29658
rect 532234 29338 532266 29574
rect 532502 29338 532586 29574
rect 532822 29338 532854 29574
rect 532234 -7066 532854 29338
rect 532234 -7302 532266 -7066
rect 532502 -7302 532586 -7066
rect 532822 -7302 532854 -7066
rect 532234 -7386 532854 -7302
rect 532234 -7622 532266 -7386
rect 532502 -7622 532586 -7386
rect 532822 -7622 532854 -7386
rect 532234 -7654 532854 -7622
rect 542194 704838 542814 711590
rect 542194 704602 542226 704838
rect 542462 704602 542546 704838
rect 542782 704602 542814 704838
rect 542194 704518 542814 704602
rect 542194 704282 542226 704518
rect 542462 704282 542546 704518
rect 542782 704282 542814 704518
rect 542194 687854 542814 704282
rect 542194 687618 542226 687854
rect 542462 687618 542546 687854
rect 542782 687618 542814 687854
rect 542194 687534 542814 687618
rect 542194 687298 542226 687534
rect 542462 687298 542546 687534
rect 542782 687298 542814 687534
rect 542194 651854 542814 687298
rect 542194 651618 542226 651854
rect 542462 651618 542546 651854
rect 542782 651618 542814 651854
rect 542194 651534 542814 651618
rect 542194 651298 542226 651534
rect 542462 651298 542546 651534
rect 542782 651298 542814 651534
rect 542194 615854 542814 651298
rect 542194 615618 542226 615854
rect 542462 615618 542546 615854
rect 542782 615618 542814 615854
rect 542194 615534 542814 615618
rect 542194 615298 542226 615534
rect 542462 615298 542546 615534
rect 542782 615298 542814 615534
rect 542194 579854 542814 615298
rect 542194 579618 542226 579854
rect 542462 579618 542546 579854
rect 542782 579618 542814 579854
rect 542194 579534 542814 579618
rect 542194 579298 542226 579534
rect 542462 579298 542546 579534
rect 542782 579298 542814 579534
rect 542194 543854 542814 579298
rect 542194 543618 542226 543854
rect 542462 543618 542546 543854
rect 542782 543618 542814 543854
rect 542194 543534 542814 543618
rect 542194 543298 542226 543534
rect 542462 543298 542546 543534
rect 542782 543298 542814 543534
rect 542194 507854 542814 543298
rect 542194 507618 542226 507854
rect 542462 507618 542546 507854
rect 542782 507618 542814 507854
rect 542194 507534 542814 507618
rect 542194 507298 542226 507534
rect 542462 507298 542546 507534
rect 542782 507298 542814 507534
rect 542194 471854 542814 507298
rect 542194 471618 542226 471854
rect 542462 471618 542546 471854
rect 542782 471618 542814 471854
rect 542194 471534 542814 471618
rect 542194 471298 542226 471534
rect 542462 471298 542546 471534
rect 542782 471298 542814 471534
rect 542194 435854 542814 471298
rect 542194 435618 542226 435854
rect 542462 435618 542546 435854
rect 542782 435618 542814 435854
rect 542194 435534 542814 435618
rect 542194 435298 542226 435534
rect 542462 435298 542546 435534
rect 542782 435298 542814 435534
rect 542194 399854 542814 435298
rect 542194 399618 542226 399854
rect 542462 399618 542546 399854
rect 542782 399618 542814 399854
rect 542194 399534 542814 399618
rect 542194 399298 542226 399534
rect 542462 399298 542546 399534
rect 542782 399298 542814 399534
rect 542194 363854 542814 399298
rect 542194 363618 542226 363854
rect 542462 363618 542546 363854
rect 542782 363618 542814 363854
rect 542194 363534 542814 363618
rect 542194 363298 542226 363534
rect 542462 363298 542546 363534
rect 542782 363298 542814 363534
rect 542194 327854 542814 363298
rect 542194 327618 542226 327854
rect 542462 327618 542546 327854
rect 542782 327618 542814 327854
rect 542194 327534 542814 327618
rect 542194 327298 542226 327534
rect 542462 327298 542546 327534
rect 542782 327298 542814 327534
rect 542194 291854 542814 327298
rect 542194 291618 542226 291854
rect 542462 291618 542546 291854
rect 542782 291618 542814 291854
rect 542194 291534 542814 291618
rect 542194 291298 542226 291534
rect 542462 291298 542546 291534
rect 542782 291298 542814 291534
rect 542194 255854 542814 291298
rect 542194 255618 542226 255854
rect 542462 255618 542546 255854
rect 542782 255618 542814 255854
rect 542194 255534 542814 255618
rect 542194 255298 542226 255534
rect 542462 255298 542546 255534
rect 542782 255298 542814 255534
rect 542194 219854 542814 255298
rect 542194 219618 542226 219854
rect 542462 219618 542546 219854
rect 542782 219618 542814 219854
rect 542194 219534 542814 219618
rect 542194 219298 542226 219534
rect 542462 219298 542546 219534
rect 542782 219298 542814 219534
rect 542194 183854 542814 219298
rect 542194 183618 542226 183854
rect 542462 183618 542546 183854
rect 542782 183618 542814 183854
rect 542194 183534 542814 183618
rect 542194 183298 542226 183534
rect 542462 183298 542546 183534
rect 542782 183298 542814 183534
rect 542194 147854 542814 183298
rect 542194 147618 542226 147854
rect 542462 147618 542546 147854
rect 542782 147618 542814 147854
rect 542194 147534 542814 147618
rect 542194 147298 542226 147534
rect 542462 147298 542546 147534
rect 542782 147298 542814 147534
rect 542194 111854 542814 147298
rect 542194 111618 542226 111854
rect 542462 111618 542546 111854
rect 542782 111618 542814 111854
rect 542194 111534 542814 111618
rect 542194 111298 542226 111534
rect 542462 111298 542546 111534
rect 542782 111298 542814 111534
rect 542194 75854 542814 111298
rect 542194 75618 542226 75854
rect 542462 75618 542546 75854
rect 542782 75618 542814 75854
rect 542194 75534 542814 75618
rect 542194 75298 542226 75534
rect 542462 75298 542546 75534
rect 542782 75298 542814 75534
rect 542194 39854 542814 75298
rect 542194 39618 542226 39854
rect 542462 39618 542546 39854
rect 542782 39618 542814 39854
rect 542194 39534 542814 39618
rect 542194 39298 542226 39534
rect 542462 39298 542546 39534
rect 542782 39298 542814 39534
rect 542194 3854 542814 39298
rect 542194 3618 542226 3854
rect 542462 3618 542546 3854
rect 542782 3618 542814 3854
rect 542194 3534 542814 3618
rect 542194 3298 542226 3534
rect 542462 3298 542546 3534
rect 542782 3298 542814 3534
rect 542194 -346 542814 3298
rect 542194 -582 542226 -346
rect 542462 -582 542546 -346
rect 542782 -582 542814 -346
rect 542194 -666 542814 -582
rect 542194 -902 542226 -666
rect 542462 -902 542546 -666
rect 542782 -902 542814 -666
rect 542194 -7654 542814 -902
rect 545914 705798 546534 711590
rect 545914 705562 545946 705798
rect 546182 705562 546266 705798
rect 546502 705562 546534 705798
rect 545914 705478 546534 705562
rect 545914 705242 545946 705478
rect 546182 705242 546266 705478
rect 546502 705242 546534 705478
rect 545914 691574 546534 705242
rect 545914 691338 545946 691574
rect 546182 691338 546266 691574
rect 546502 691338 546534 691574
rect 545914 691254 546534 691338
rect 545914 691018 545946 691254
rect 546182 691018 546266 691254
rect 546502 691018 546534 691254
rect 545914 655574 546534 691018
rect 545914 655338 545946 655574
rect 546182 655338 546266 655574
rect 546502 655338 546534 655574
rect 545914 655254 546534 655338
rect 545914 655018 545946 655254
rect 546182 655018 546266 655254
rect 546502 655018 546534 655254
rect 545914 619574 546534 655018
rect 545914 619338 545946 619574
rect 546182 619338 546266 619574
rect 546502 619338 546534 619574
rect 545914 619254 546534 619338
rect 545914 619018 545946 619254
rect 546182 619018 546266 619254
rect 546502 619018 546534 619254
rect 545914 583574 546534 619018
rect 545914 583338 545946 583574
rect 546182 583338 546266 583574
rect 546502 583338 546534 583574
rect 545914 583254 546534 583338
rect 545914 583018 545946 583254
rect 546182 583018 546266 583254
rect 546502 583018 546534 583254
rect 545914 547574 546534 583018
rect 545914 547338 545946 547574
rect 546182 547338 546266 547574
rect 546502 547338 546534 547574
rect 545914 547254 546534 547338
rect 545914 547018 545946 547254
rect 546182 547018 546266 547254
rect 546502 547018 546534 547254
rect 545914 511574 546534 547018
rect 545914 511338 545946 511574
rect 546182 511338 546266 511574
rect 546502 511338 546534 511574
rect 545914 511254 546534 511338
rect 545914 511018 545946 511254
rect 546182 511018 546266 511254
rect 546502 511018 546534 511254
rect 545914 475574 546534 511018
rect 545914 475338 545946 475574
rect 546182 475338 546266 475574
rect 546502 475338 546534 475574
rect 545914 475254 546534 475338
rect 545914 475018 545946 475254
rect 546182 475018 546266 475254
rect 546502 475018 546534 475254
rect 545914 439574 546534 475018
rect 545914 439338 545946 439574
rect 546182 439338 546266 439574
rect 546502 439338 546534 439574
rect 545914 439254 546534 439338
rect 545914 439018 545946 439254
rect 546182 439018 546266 439254
rect 546502 439018 546534 439254
rect 545914 403574 546534 439018
rect 545914 403338 545946 403574
rect 546182 403338 546266 403574
rect 546502 403338 546534 403574
rect 545914 403254 546534 403338
rect 545914 403018 545946 403254
rect 546182 403018 546266 403254
rect 546502 403018 546534 403254
rect 545914 367574 546534 403018
rect 545914 367338 545946 367574
rect 546182 367338 546266 367574
rect 546502 367338 546534 367574
rect 545914 367254 546534 367338
rect 545914 367018 545946 367254
rect 546182 367018 546266 367254
rect 546502 367018 546534 367254
rect 545914 331574 546534 367018
rect 545914 331338 545946 331574
rect 546182 331338 546266 331574
rect 546502 331338 546534 331574
rect 545914 331254 546534 331338
rect 545914 331018 545946 331254
rect 546182 331018 546266 331254
rect 546502 331018 546534 331254
rect 545914 295574 546534 331018
rect 545914 295338 545946 295574
rect 546182 295338 546266 295574
rect 546502 295338 546534 295574
rect 545914 295254 546534 295338
rect 545914 295018 545946 295254
rect 546182 295018 546266 295254
rect 546502 295018 546534 295254
rect 545914 259574 546534 295018
rect 545914 259338 545946 259574
rect 546182 259338 546266 259574
rect 546502 259338 546534 259574
rect 545914 259254 546534 259338
rect 545914 259018 545946 259254
rect 546182 259018 546266 259254
rect 546502 259018 546534 259254
rect 545914 223574 546534 259018
rect 545914 223338 545946 223574
rect 546182 223338 546266 223574
rect 546502 223338 546534 223574
rect 545914 223254 546534 223338
rect 545914 223018 545946 223254
rect 546182 223018 546266 223254
rect 546502 223018 546534 223254
rect 545914 187574 546534 223018
rect 545914 187338 545946 187574
rect 546182 187338 546266 187574
rect 546502 187338 546534 187574
rect 545914 187254 546534 187338
rect 545914 187018 545946 187254
rect 546182 187018 546266 187254
rect 546502 187018 546534 187254
rect 545914 151574 546534 187018
rect 545914 151338 545946 151574
rect 546182 151338 546266 151574
rect 546502 151338 546534 151574
rect 545914 151254 546534 151338
rect 545914 151018 545946 151254
rect 546182 151018 546266 151254
rect 546502 151018 546534 151254
rect 545914 115574 546534 151018
rect 545914 115338 545946 115574
rect 546182 115338 546266 115574
rect 546502 115338 546534 115574
rect 545914 115254 546534 115338
rect 545914 115018 545946 115254
rect 546182 115018 546266 115254
rect 546502 115018 546534 115254
rect 545914 79574 546534 115018
rect 545914 79338 545946 79574
rect 546182 79338 546266 79574
rect 546502 79338 546534 79574
rect 545914 79254 546534 79338
rect 545914 79018 545946 79254
rect 546182 79018 546266 79254
rect 546502 79018 546534 79254
rect 545914 43574 546534 79018
rect 545914 43338 545946 43574
rect 546182 43338 546266 43574
rect 546502 43338 546534 43574
rect 545914 43254 546534 43338
rect 545914 43018 545946 43254
rect 546182 43018 546266 43254
rect 546502 43018 546534 43254
rect 545914 7574 546534 43018
rect 545914 7338 545946 7574
rect 546182 7338 546266 7574
rect 546502 7338 546534 7574
rect 545914 7254 546534 7338
rect 545914 7018 545946 7254
rect 546182 7018 546266 7254
rect 546502 7018 546534 7254
rect 545914 -1306 546534 7018
rect 545914 -1542 545946 -1306
rect 546182 -1542 546266 -1306
rect 546502 -1542 546534 -1306
rect 545914 -1626 546534 -1542
rect 545914 -1862 545946 -1626
rect 546182 -1862 546266 -1626
rect 546502 -1862 546534 -1626
rect 545914 -7654 546534 -1862
rect 549634 706758 550254 711590
rect 549634 706522 549666 706758
rect 549902 706522 549986 706758
rect 550222 706522 550254 706758
rect 549634 706438 550254 706522
rect 549634 706202 549666 706438
rect 549902 706202 549986 706438
rect 550222 706202 550254 706438
rect 549634 695294 550254 706202
rect 549634 695058 549666 695294
rect 549902 695058 549986 695294
rect 550222 695058 550254 695294
rect 549634 694974 550254 695058
rect 549634 694738 549666 694974
rect 549902 694738 549986 694974
rect 550222 694738 550254 694974
rect 549634 659294 550254 694738
rect 549634 659058 549666 659294
rect 549902 659058 549986 659294
rect 550222 659058 550254 659294
rect 549634 658974 550254 659058
rect 549634 658738 549666 658974
rect 549902 658738 549986 658974
rect 550222 658738 550254 658974
rect 549634 623294 550254 658738
rect 549634 623058 549666 623294
rect 549902 623058 549986 623294
rect 550222 623058 550254 623294
rect 549634 622974 550254 623058
rect 549634 622738 549666 622974
rect 549902 622738 549986 622974
rect 550222 622738 550254 622974
rect 549634 587294 550254 622738
rect 549634 587058 549666 587294
rect 549902 587058 549986 587294
rect 550222 587058 550254 587294
rect 549634 586974 550254 587058
rect 549634 586738 549666 586974
rect 549902 586738 549986 586974
rect 550222 586738 550254 586974
rect 549634 551294 550254 586738
rect 549634 551058 549666 551294
rect 549902 551058 549986 551294
rect 550222 551058 550254 551294
rect 549634 550974 550254 551058
rect 549634 550738 549666 550974
rect 549902 550738 549986 550974
rect 550222 550738 550254 550974
rect 549634 515294 550254 550738
rect 549634 515058 549666 515294
rect 549902 515058 549986 515294
rect 550222 515058 550254 515294
rect 549634 514974 550254 515058
rect 549634 514738 549666 514974
rect 549902 514738 549986 514974
rect 550222 514738 550254 514974
rect 549634 479294 550254 514738
rect 549634 479058 549666 479294
rect 549902 479058 549986 479294
rect 550222 479058 550254 479294
rect 549634 478974 550254 479058
rect 549634 478738 549666 478974
rect 549902 478738 549986 478974
rect 550222 478738 550254 478974
rect 549634 443294 550254 478738
rect 549634 443058 549666 443294
rect 549902 443058 549986 443294
rect 550222 443058 550254 443294
rect 549634 442974 550254 443058
rect 549634 442738 549666 442974
rect 549902 442738 549986 442974
rect 550222 442738 550254 442974
rect 549634 407294 550254 442738
rect 549634 407058 549666 407294
rect 549902 407058 549986 407294
rect 550222 407058 550254 407294
rect 549634 406974 550254 407058
rect 549634 406738 549666 406974
rect 549902 406738 549986 406974
rect 550222 406738 550254 406974
rect 549634 371294 550254 406738
rect 549634 371058 549666 371294
rect 549902 371058 549986 371294
rect 550222 371058 550254 371294
rect 549634 370974 550254 371058
rect 549634 370738 549666 370974
rect 549902 370738 549986 370974
rect 550222 370738 550254 370974
rect 549634 335294 550254 370738
rect 549634 335058 549666 335294
rect 549902 335058 549986 335294
rect 550222 335058 550254 335294
rect 549634 334974 550254 335058
rect 549634 334738 549666 334974
rect 549902 334738 549986 334974
rect 550222 334738 550254 334974
rect 549634 299294 550254 334738
rect 549634 299058 549666 299294
rect 549902 299058 549986 299294
rect 550222 299058 550254 299294
rect 549634 298974 550254 299058
rect 549634 298738 549666 298974
rect 549902 298738 549986 298974
rect 550222 298738 550254 298974
rect 549634 263294 550254 298738
rect 549634 263058 549666 263294
rect 549902 263058 549986 263294
rect 550222 263058 550254 263294
rect 549634 262974 550254 263058
rect 549634 262738 549666 262974
rect 549902 262738 549986 262974
rect 550222 262738 550254 262974
rect 549634 227294 550254 262738
rect 549634 227058 549666 227294
rect 549902 227058 549986 227294
rect 550222 227058 550254 227294
rect 549634 226974 550254 227058
rect 549634 226738 549666 226974
rect 549902 226738 549986 226974
rect 550222 226738 550254 226974
rect 549634 191294 550254 226738
rect 549634 191058 549666 191294
rect 549902 191058 549986 191294
rect 550222 191058 550254 191294
rect 549634 190974 550254 191058
rect 549634 190738 549666 190974
rect 549902 190738 549986 190974
rect 550222 190738 550254 190974
rect 549634 155294 550254 190738
rect 549634 155058 549666 155294
rect 549902 155058 549986 155294
rect 550222 155058 550254 155294
rect 549634 154974 550254 155058
rect 549634 154738 549666 154974
rect 549902 154738 549986 154974
rect 550222 154738 550254 154974
rect 549634 119294 550254 154738
rect 549634 119058 549666 119294
rect 549902 119058 549986 119294
rect 550222 119058 550254 119294
rect 549634 118974 550254 119058
rect 549634 118738 549666 118974
rect 549902 118738 549986 118974
rect 550222 118738 550254 118974
rect 549634 83294 550254 118738
rect 549634 83058 549666 83294
rect 549902 83058 549986 83294
rect 550222 83058 550254 83294
rect 549634 82974 550254 83058
rect 549634 82738 549666 82974
rect 549902 82738 549986 82974
rect 550222 82738 550254 82974
rect 549634 47294 550254 82738
rect 549634 47058 549666 47294
rect 549902 47058 549986 47294
rect 550222 47058 550254 47294
rect 549634 46974 550254 47058
rect 549634 46738 549666 46974
rect 549902 46738 549986 46974
rect 550222 46738 550254 46974
rect 549634 11294 550254 46738
rect 549634 11058 549666 11294
rect 549902 11058 549986 11294
rect 550222 11058 550254 11294
rect 549634 10974 550254 11058
rect 549634 10738 549666 10974
rect 549902 10738 549986 10974
rect 550222 10738 550254 10974
rect 549634 -2266 550254 10738
rect 549634 -2502 549666 -2266
rect 549902 -2502 549986 -2266
rect 550222 -2502 550254 -2266
rect 549634 -2586 550254 -2502
rect 549634 -2822 549666 -2586
rect 549902 -2822 549986 -2586
rect 550222 -2822 550254 -2586
rect 549634 -7654 550254 -2822
rect 553354 707718 553974 711590
rect 553354 707482 553386 707718
rect 553622 707482 553706 707718
rect 553942 707482 553974 707718
rect 553354 707398 553974 707482
rect 553354 707162 553386 707398
rect 553622 707162 553706 707398
rect 553942 707162 553974 707398
rect 553354 699014 553974 707162
rect 553354 698778 553386 699014
rect 553622 698778 553706 699014
rect 553942 698778 553974 699014
rect 553354 698694 553974 698778
rect 553354 698458 553386 698694
rect 553622 698458 553706 698694
rect 553942 698458 553974 698694
rect 553354 663014 553974 698458
rect 553354 662778 553386 663014
rect 553622 662778 553706 663014
rect 553942 662778 553974 663014
rect 553354 662694 553974 662778
rect 553354 662458 553386 662694
rect 553622 662458 553706 662694
rect 553942 662458 553974 662694
rect 553354 627014 553974 662458
rect 553354 626778 553386 627014
rect 553622 626778 553706 627014
rect 553942 626778 553974 627014
rect 553354 626694 553974 626778
rect 553354 626458 553386 626694
rect 553622 626458 553706 626694
rect 553942 626458 553974 626694
rect 553354 591014 553974 626458
rect 553354 590778 553386 591014
rect 553622 590778 553706 591014
rect 553942 590778 553974 591014
rect 553354 590694 553974 590778
rect 553354 590458 553386 590694
rect 553622 590458 553706 590694
rect 553942 590458 553974 590694
rect 553354 555014 553974 590458
rect 553354 554778 553386 555014
rect 553622 554778 553706 555014
rect 553942 554778 553974 555014
rect 553354 554694 553974 554778
rect 553354 554458 553386 554694
rect 553622 554458 553706 554694
rect 553942 554458 553974 554694
rect 553354 519014 553974 554458
rect 553354 518778 553386 519014
rect 553622 518778 553706 519014
rect 553942 518778 553974 519014
rect 553354 518694 553974 518778
rect 553354 518458 553386 518694
rect 553622 518458 553706 518694
rect 553942 518458 553974 518694
rect 553354 483014 553974 518458
rect 553354 482778 553386 483014
rect 553622 482778 553706 483014
rect 553942 482778 553974 483014
rect 553354 482694 553974 482778
rect 553354 482458 553386 482694
rect 553622 482458 553706 482694
rect 553942 482458 553974 482694
rect 553354 447014 553974 482458
rect 553354 446778 553386 447014
rect 553622 446778 553706 447014
rect 553942 446778 553974 447014
rect 553354 446694 553974 446778
rect 553354 446458 553386 446694
rect 553622 446458 553706 446694
rect 553942 446458 553974 446694
rect 553354 411014 553974 446458
rect 553354 410778 553386 411014
rect 553622 410778 553706 411014
rect 553942 410778 553974 411014
rect 553354 410694 553974 410778
rect 553354 410458 553386 410694
rect 553622 410458 553706 410694
rect 553942 410458 553974 410694
rect 553354 375014 553974 410458
rect 553354 374778 553386 375014
rect 553622 374778 553706 375014
rect 553942 374778 553974 375014
rect 553354 374694 553974 374778
rect 553354 374458 553386 374694
rect 553622 374458 553706 374694
rect 553942 374458 553974 374694
rect 553354 339014 553974 374458
rect 553354 338778 553386 339014
rect 553622 338778 553706 339014
rect 553942 338778 553974 339014
rect 553354 338694 553974 338778
rect 553354 338458 553386 338694
rect 553622 338458 553706 338694
rect 553942 338458 553974 338694
rect 553354 303014 553974 338458
rect 553354 302778 553386 303014
rect 553622 302778 553706 303014
rect 553942 302778 553974 303014
rect 553354 302694 553974 302778
rect 553354 302458 553386 302694
rect 553622 302458 553706 302694
rect 553942 302458 553974 302694
rect 553354 267014 553974 302458
rect 553354 266778 553386 267014
rect 553622 266778 553706 267014
rect 553942 266778 553974 267014
rect 553354 266694 553974 266778
rect 553354 266458 553386 266694
rect 553622 266458 553706 266694
rect 553942 266458 553974 266694
rect 553354 231014 553974 266458
rect 553354 230778 553386 231014
rect 553622 230778 553706 231014
rect 553942 230778 553974 231014
rect 553354 230694 553974 230778
rect 553354 230458 553386 230694
rect 553622 230458 553706 230694
rect 553942 230458 553974 230694
rect 553354 195014 553974 230458
rect 553354 194778 553386 195014
rect 553622 194778 553706 195014
rect 553942 194778 553974 195014
rect 553354 194694 553974 194778
rect 553354 194458 553386 194694
rect 553622 194458 553706 194694
rect 553942 194458 553974 194694
rect 553354 159014 553974 194458
rect 553354 158778 553386 159014
rect 553622 158778 553706 159014
rect 553942 158778 553974 159014
rect 553354 158694 553974 158778
rect 553354 158458 553386 158694
rect 553622 158458 553706 158694
rect 553942 158458 553974 158694
rect 553354 123014 553974 158458
rect 553354 122778 553386 123014
rect 553622 122778 553706 123014
rect 553942 122778 553974 123014
rect 553354 122694 553974 122778
rect 553354 122458 553386 122694
rect 553622 122458 553706 122694
rect 553942 122458 553974 122694
rect 553354 87014 553974 122458
rect 553354 86778 553386 87014
rect 553622 86778 553706 87014
rect 553942 86778 553974 87014
rect 553354 86694 553974 86778
rect 553354 86458 553386 86694
rect 553622 86458 553706 86694
rect 553942 86458 553974 86694
rect 553354 51014 553974 86458
rect 553354 50778 553386 51014
rect 553622 50778 553706 51014
rect 553942 50778 553974 51014
rect 553354 50694 553974 50778
rect 553354 50458 553386 50694
rect 553622 50458 553706 50694
rect 553942 50458 553974 50694
rect 553354 15014 553974 50458
rect 553354 14778 553386 15014
rect 553622 14778 553706 15014
rect 553942 14778 553974 15014
rect 553354 14694 553974 14778
rect 553354 14458 553386 14694
rect 553622 14458 553706 14694
rect 553942 14458 553974 14694
rect 553354 -3226 553974 14458
rect 553354 -3462 553386 -3226
rect 553622 -3462 553706 -3226
rect 553942 -3462 553974 -3226
rect 553354 -3546 553974 -3462
rect 553354 -3782 553386 -3546
rect 553622 -3782 553706 -3546
rect 553942 -3782 553974 -3546
rect 553354 -7654 553974 -3782
rect 557074 708678 557694 711590
rect 557074 708442 557106 708678
rect 557342 708442 557426 708678
rect 557662 708442 557694 708678
rect 557074 708358 557694 708442
rect 557074 708122 557106 708358
rect 557342 708122 557426 708358
rect 557662 708122 557694 708358
rect 557074 666734 557694 708122
rect 557074 666498 557106 666734
rect 557342 666498 557426 666734
rect 557662 666498 557694 666734
rect 557074 666414 557694 666498
rect 557074 666178 557106 666414
rect 557342 666178 557426 666414
rect 557662 666178 557694 666414
rect 557074 630734 557694 666178
rect 557074 630498 557106 630734
rect 557342 630498 557426 630734
rect 557662 630498 557694 630734
rect 557074 630414 557694 630498
rect 557074 630178 557106 630414
rect 557342 630178 557426 630414
rect 557662 630178 557694 630414
rect 557074 594734 557694 630178
rect 557074 594498 557106 594734
rect 557342 594498 557426 594734
rect 557662 594498 557694 594734
rect 557074 594414 557694 594498
rect 557074 594178 557106 594414
rect 557342 594178 557426 594414
rect 557662 594178 557694 594414
rect 557074 558734 557694 594178
rect 557074 558498 557106 558734
rect 557342 558498 557426 558734
rect 557662 558498 557694 558734
rect 557074 558414 557694 558498
rect 557074 558178 557106 558414
rect 557342 558178 557426 558414
rect 557662 558178 557694 558414
rect 557074 522734 557694 558178
rect 557074 522498 557106 522734
rect 557342 522498 557426 522734
rect 557662 522498 557694 522734
rect 557074 522414 557694 522498
rect 557074 522178 557106 522414
rect 557342 522178 557426 522414
rect 557662 522178 557694 522414
rect 557074 486734 557694 522178
rect 557074 486498 557106 486734
rect 557342 486498 557426 486734
rect 557662 486498 557694 486734
rect 557074 486414 557694 486498
rect 557074 486178 557106 486414
rect 557342 486178 557426 486414
rect 557662 486178 557694 486414
rect 557074 450734 557694 486178
rect 557074 450498 557106 450734
rect 557342 450498 557426 450734
rect 557662 450498 557694 450734
rect 557074 450414 557694 450498
rect 557074 450178 557106 450414
rect 557342 450178 557426 450414
rect 557662 450178 557694 450414
rect 557074 414734 557694 450178
rect 557074 414498 557106 414734
rect 557342 414498 557426 414734
rect 557662 414498 557694 414734
rect 557074 414414 557694 414498
rect 557074 414178 557106 414414
rect 557342 414178 557426 414414
rect 557662 414178 557694 414414
rect 557074 378734 557694 414178
rect 557074 378498 557106 378734
rect 557342 378498 557426 378734
rect 557662 378498 557694 378734
rect 557074 378414 557694 378498
rect 557074 378178 557106 378414
rect 557342 378178 557426 378414
rect 557662 378178 557694 378414
rect 557074 342734 557694 378178
rect 557074 342498 557106 342734
rect 557342 342498 557426 342734
rect 557662 342498 557694 342734
rect 557074 342414 557694 342498
rect 557074 342178 557106 342414
rect 557342 342178 557426 342414
rect 557662 342178 557694 342414
rect 557074 306734 557694 342178
rect 557074 306498 557106 306734
rect 557342 306498 557426 306734
rect 557662 306498 557694 306734
rect 557074 306414 557694 306498
rect 557074 306178 557106 306414
rect 557342 306178 557426 306414
rect 557662 306178 557694 306414
rect 557074 270734 557694 306178
rect 557074 270498 557106 270734
rect 557342 270498 557426 270734
rect 557662 270498 557694 270734
rect 557074 270414 557694 270498
rect 557074 270178 557106 270414
rect 557342 270178 557426 270414
rect 557662 270178 557694 270414
rect 557074 234734 557694 270178
rect 557074 234498 557106 234734
rect 557342 234498 557426 234734
rect 557662 234498 557694 234734
rect 557074 234414 557694 234498
rect 557074 234178 557106 234414
rect 557342 234178 557426 234414
rect 557662 234178 557694 234414
rect 557074 198734 557694 234178
rect 557074 198498 557106 198734
rect 557342 198498 557426 198734
rect 557662 198498 557694 198734
rect 557074 198414 557694 198498
rect 557074 198178 557106 198414
rect 557342 198178 557426 198414
rect 557662 198178 557694 198414
rect 557074 162734 557694 198178
rect 557074 162498 557106 162734
rect 557342 162498 557426 162734
rect 557662 162498 557694 162734
rect 557074 162414 557694 162498
rect 557074 162178 557106 162414
rect 557342 162178 557426 162414
rect 557662 162178 557694 162414
rect 557074 126734 557694 162178
rect 557074 126498 557106 126734
rect 557342 126498 557426 126734
rect 557662 126498 557694 126734
rect 557074 126414 557694 126498
rect 557074 126178 557106 126414
rect 557342 126178 557426 126414
rect 557662 126178 557694 126414
rect 557074 90734 557694 126178
rect 557074 90498 557106 90734
rect 557342 90498 557426 90734
rect 557662 90498 557694 90734
rect 557074 90414 557694 90498
rect 557074 90178 557106 90414
rect 557342 90178 557426 90414
rect 557662 90178 557694 90414
rect 557074 54734 557694 90178
rect 557074 54498 557106 54734
rect 557342 54498 557426 54734
rect 557662 54498 557694 54734
rect 557074 54414 557694 54498
rect 557074 54178 557106 54414
rect 557342 54178 557426 54414
rect 557662 54178 557694 54414
rect 557074 18734 557694 54178
rect 557074 18498 557106 18734
rect 557342 18498 557426 18734
rect 557662 18498 557694 18734
rect 557074 18414 557694 18498
rect 557074 18178 557106 18414
rect 557342 18178 557426 18414
rect 557662 18178 557694 18414
rect 557074 -4186 557694 18178
rect 557074 -4422 557106 -4186
rect 557342 -4422 557426 -4186
rect 557662 -4422 557694 -4186
rect 557074 -4506 557694 -4422
rect 557074 -4742 557106 -4506
rect 557342 -4742 557426 -4506
rect 557662 -4742 557694 -4506
rect 557074 -7654 557694 -4742
rect 560794 709638 561414 711590
rect 560794 709402 560826 709638
rect 561062 709402 561146 709638
rect 561382 709402 561414 709638
rect 560794 709318 561414 709402
rect 560794 709082 560826 709318
rect 561062 709082 561146 709318
rect 561382 709082 561414 709318
rect 560794 670454 561414 709082
rect 560794 670218 560826 670454
rect 561062 670218 561146 670454
rect 561382 670218 561414 670454
rect 560794 670134 561414 670218
rect 560794 669898 560826 670134
rect 561062 669898 561146 670134
rect 561382 669898 561414 670134
rect 560794 634454 561414 669898
rect 560794 634218 560826 634454
rect 561062 634218 561146 634454
rect 561382 634218 561414 634454
rect 560794 634134 561414 634218
rect 560794 633898 560826 634134
rect 561062 633898 561146 634134
rect 561382 633898 561414 634134
rect 560794 598454 561414 633898
rect 560794 598218 560826 598454
rect 561062 598218 561146 598454
rect 561382 598218 561414 598454
rect 560794 598134 561414 598218
rect 560794 597898 560826 598134
rect 561062 597898 561146 598134
rect 561382 597898 561414 598134
rect 560794 562454 561414 597898
rect 560794 562218 560826 562454
rect 561062 562218 561146 562454
rect 561382 562218 561414 562454
rect 560794 562134 561414 562218
rect 560794 561898 560826 562134
rect 561062 561898 561146 562134
rect 561382 561898 561414 562134
rect 560794 526454 561414 561898
rect 560794 526218 560826 526454
rect 561062 526218 561146 526454
rect 561382 526218 561414 526454
rect 560794 526134 561414 526218
rect 560794 525898 560826 526134
rect 561062 525898 561146 526134
rect 561382 525898 561414 526134
rect 560794 490454 561414 525898
rect 560794 490218 560826 490454
rect 561062 490218 561146 490454
rect 561382 490218 561414 490454
rect 560794 490134 561414 490218
rect 560794 489898 560826 490134
rect 561062 489898 561146 490134
rect 561382 489898 561414 490134
rect 560794 454454 561414 489898
rect 560794 454218 560826 454454
rect 561062 454218 561146 454454
rect 561382 454218 561414 454454
rect 560794 454134 561414 454218
rect 560794 453898 560826 454134
rect 561062 453898 561146 454134
rect 561382 453898 561414 454134
rect 560794 418454 561414 453898
rect 560794 418218 560826 418454
rect 561062 418218 561146 418454
rect 561382 418218 561414 418454
rect 560794 418134 561414 418218
rect 560794 417898 560826 418134
rect 561062 417898 561146 418134
rect 561382 417898 561414 418134
rect 560794 382454 561414 417898
rect 560794 382218 560826 382454
rect 561062 382218 561146 382454
rect 561382 382218 561414 382454
rect 560794 382134 561414 382218
rect 560794 381898 560826 382134
rect 561062 381898 561146 382134
rect 561382 381898 561414 382134
rect 560794 346454 561414 381898
rect 560794 346218 560826 346454
rect 561062 346218 561146 346454
rect 561382 346218 561414 346454
rect 560794 346134 561414 346218
rect 560794 345898 560826 346134
rect 561062 345898 561146 346134
rect 561382 345898 561414 346134
rect 560794 310454 561414 345898
rect 560794 310218 560826 310454
rect 561062 310218 561146 310454
rect 561382 310218 561414 310454
rect 560794 310134 561414 310218
rect 560794 309898 560826 310134
rect 561062 309898 561146 310134
rect 561382 309898 561414 310134
rect 560794 274454 561414 309898
rect 560794 274218 560826 274454
rect 561062 274218 561146 274454
rect 561382 274218 561414 274454
rect 560794 274134 561414 274218
rect 560794 273898 560826 274134
rect 561062 273898 561146 274134
rect 561382 273898 561414 274134
rect 560794 238454 561414 273898
rect 560794 238218 560826 238454
rect 561062 238218 561146 238454
rect 561382 238218 561414 238454
rect 560794 238134 561414 238218
rect 560794 237898 560826 238134
rect 561062 237898 561146 238134
rect 561382 237898 561414 238134
rect 560794 202454 561414 237898
rect 560794 202218 560826 202454
rect 561062 202218 561146 202454
rect 561382 202218 561414 202454
rect 560794 202134 561414 202218
rect 560794 201898 560826 202134
rect 561062 201898 561146 202134
rect 561382 201898 561414 202134
rect 560794 166454 561414 201898
rect 560794 166218 560826 166454
rect 561062 166218 561146 166454
rect 561382 166218 561414 166454
rect 560794 166134 561414 166218
rect 560794 165898 560826 166134
rect 561062 165898 561146 166134
rect 561382 165898 561414 166134
rect 560794 130454 561414 165898
rect 560794 130218 560826 130454
rect 561062 130218 561146 130454
rect 561382 130218 561414 130454
rect 560794 130134 561414 130218
rect 560794 129898 560826 130134
rect 561062 129898 561146 130134
rect 561382 129898 561414 130134
rect 560794 94454 561414 129898
rect 560794 94218 560826 94454
rect 561062 94218 561146 94454
rect 561382 94218 561414 94454
rect 560794 94134 561414 94218
rect 560794 93898 560826 94134
rect 561062 93898 561146 94134
rect 561382 93898 561414 94134
rect 560794 58454 561414 93898
rect 560794 58218 560826 58454
rect 561062 58218 561146 58454
rect 561382 58218 561414 58454
rect 560794 58134 561414 58218
rect 560794 57898 560826 58134
rect 561062 57898 561146 58134
rect 561382 57898 561414 58134
rect 560794 22454 561414 57898
rect 560794 22218 560826 22454
rect 561062 22218 561146 22454
rect 561382 22218 561414 22454
rect 560794 22134 561414 22218
rect 560794 21898 560826 22134
rect 561062 21898 561146 22134
rect 561382 21898 561414 22134
rect 560794 -5146 561414 21898
rect 560794 -5382 560826 -5146
rect 561062 -5382 561146 -5146
rect 561382 -5382 561414 -5146
rect 560794 -5466 561414 -5382
rect 560794 -5702 560826 -5466
rect 561062 -5702 561146 -5466
rect 561382 -5702 561414 -5466
rect 560794 -7654 561414 -5702
rect 564514 710598 565134 711590
rect 564514 710362 564546 710598
rect 564782 710362 564866 710598
rect 565102 710362 565134 710598
rect 564514 710278 565134 710362
rect 564514 710042 564546 710278
rect 564782 710042 564866 710278
rect 565102 710042 565134 710278
rect 564514 674174 565134 710042
rect 564514 673938 564546 674174
rect 564782 673938 564866 674174
rect 565102 673938 565134 674174
rect 564514 673854 565134 673938
rect 564514 673618 564546 673854
rect 564782 673618 564866 673854
rect 565102 673618 565134 673854
rect 564514 638174 565134 673618
rect 564514 637938 564546 638174
rect 564782 637938 564866 638174
rect 565102 637938 565134 638174
rect 564514 637854 565134 637938
rect 564514 637618 564546 637854
rect 564782 637618 564866 637854
rect 565102 637618 565134 637854
rect 564514 602174 565134 637618
rect 564514 601938 564546 602174
rect 564782 601938 564866 602174
rect 565102 601938 565134 602174
rect 564514 601854 565134 601938
rect 564514 601618 564546 601854
rect 564782 601618 564866 601854
rect 565102 601618 565134 601854
rect 564514 566174 565134 601618
rect 564514 565938 564546 566174
rect 564782 565938 564866 566174
rect 565102 565938 565134 566174
rect 564514 565854 565134 565938
rect 564514 565618 564546 565854
rect 564782 565618 564866 565854
rect 565102 565618 565134 565854
rect 564514 530174 565134 565618
rect 564514 529938 564546 530174
rect 564782 529938 564866 530174
rect 565102 529938 565134 530174
rect 564514 529854 565134 529938
rect 564514 529618 564546 529854
rect 564782 529618 564866 529854
rect 565102 529618 565134 529854
rect 564514 494174 565134 529618
rect 564514 493938 564546 494174
rect 564782 493938 564866 494174
rect 565102 493938 565134 494174
rect 564514 493854 565134 493938
rect 564514 493618 564546 493854
rect 564782 493618 564866 493854
rect 565102 493618 565134 493854
rect 564514 458174 565134 493618
rect 564514 457938 564546 458174
rect 564782 457938 564866 458174
rect 565102 457938 565134 458174
rect 564514 457854 565134 457938
rect 564514 457618 564546 457854
rect 564782 457618 564866 457854
rect 565102 457618 565134 457854
rect 564514 422174 565134 457618
rect 564514 421938 564546 422174
rect 564782 421938 564866 422174
rect 565102 421938 565134 422174
rect 564514 421854 565134 421938
rect 564514 421618 564546 421854
rect 564782 421618 564866 421854
rect 565102 421618 565134 421854
rect 564514 386174 565134 421618
rect 564514 385938 564546 386174
rect 564782 385938 564866 386174
rect 565102 385938 565134 386174
rect 564514 385854 565134 385938
rect 564514 385618 564546 385854
rect 564782 385618 564866 385854
rect 565102 385618 565134 385854
rect 564514 350174 565134 385618
rect 564514 349938 564546 350174
rect 564782 349938 564866 350174
rect 565102 349938 565134 350174
rect 564514 349854 565134 349938
rect 564514 349618 564546 349854
rect 564782 349618 564866 349854
rect 565102 349618 565134 349854
rect 564514 314174 565134 349618
rect 564514 313938 564546 314174
rect 564782 313938 564866 314174
rect 565102 313938 565134 314174
rect 564514 313854 565134 313938
rect 564514 313618 564546 313854
rect 564782 313618 564866 313854
rect 565102 313618 565134 313854
rect 564514 278174 565134 313618
rect 564514 277938 564546 278174
rect 564782 277938 564866 278174
rect 565102 277938 565134 278174
rect 564514 277854 565134 277938
rect 564514 277618 564546 277854
rect 564782 277618 564866 277854
rect 565102 277618 565134 277854
rect 564514 242174 565134 277618
rect 564514 241938 564546 242174
rect 564782 241938 564866 242174
rect 565102 241938 565134 242174
rect 564514 241854 565134 241938
rect 564514 241618 564546 241854
rect 564782 241618 564866 241854
rect 565102 241618 565134 241854
rect 564514 206174 565134 241618
rect 564514 205938 564546 206174
rect 564782 205938 564866 206174
rect 565102 205938 565134 206174
rect 564514 205854 565134 205938
rect 564514 205618 564546 205854
rect 564782 205618 564866 205854
rect 565102 205618 565134 205854
rect 564514 170174 565134 205618
rect 564514 169938 564546 170174
rect 564782 169938 564866 170174
rect 565102 169938 565134 170174
rect 564514 169854 565134 169938
rect 564514 169618 564546 169854
rect 564782 169618 564866 169854
rect 565102 169618 565134 169854
rect 564514 134174 565134 169618
rect 564514 133938 564546 134174
rect 564782 133938 564866 134174
rect 565102 133938 565134 134174
rect 564514 133854 565134 133938
rect 564514 133618 564546 133854
rect 564782 133618 564866 133854
rect 565102 133618 565134 133854
rect 564514 98174 565134 133618
rect 564514 97938 564546 98174
rect 564782 97938 564866 98174
rect 565102 97938 565134 98174
rect 564514 97854 565134 97938
rect 564514 97618 564546 97854
rect 564782 97618 564866 97854
rect 565102 97618 565134 97854
rect 564514 62174 565134 97618
rect 564514 61938 564546 62174
rect 564782 61938 564866 62174
rect 565102 61938 565134 62174
rect 564514 61854 565134 61938
rect 564514 61618 564546 61854
rect 564782 61618 564866 61854
rect 565102 61618 565134 61854
rect 564514 26174 565134 61618
rect 564514 25938 564546 26174
rect 564782 25938 564866 26174
rect 565102 25938 565134 26174
rect 564514 25854 565134 25938
rect 564514 25618 564546 25854
rect 564782 25618 564866 25854
rect 565102 25618 565134 25854
rect 564514 -6106 565134 25618
rect 564514 -6342 564546 -6106
rect 564782 -6342 564866 -6106
rect 565102 -6342 565134 -6106
rect 564514 -6426 565134 -6342
rect 564514 -6662 564546 -6426
rect 564782 -6662 564866 -6426
rect 565102 -6662 565134 -6426
rect 564514 -7654 565134 -6662
rect 568234 711558 568854 711590
rect 568234 711322 568266 711558
rect 568502 711322 568586 711558
rect 568822 711322 568854 711558
rect 568234 711238 568854 711322
rect 568234 711002 568266 711238
rect 568502 711002 568586 711238
rect 568822 711002 568854 711238
rect 568234 677894 568854 711002
rect 568234 677658 568266 677894
rect 568502 677658 568586 677894
rect 568822 677658 568854 677894
rect 568234 677574 568854 677658
rect 568234 677338 568266 677574
rect 568502 677338 568586 677574
rect 568822 677338 568854 677574
rect 568234 641894 568854 677338
rect 568234 641658 568266 641894
rect 568502 641658 568586 641894
rect 568822 641658 568854 641894
rect 568234 641574 568854 641658
rect 568234 641338 568266 641574
rect 568502 641338 568586 641574
rect 568822 641338 568854 641574
rect 568234 605894 568854 641338
rect 568234 605658 568266 605894
rect 568502 605658 568586 605894
rect 568822 605658 568854 605894
rect 568234 605574 568854 605658
rect 568234 605338 568266 605574
rect 568502 605338 568586 605574
rect 568822 605338 568854 605574
rect 568234 569894 568854 605338
rect 568234 569658 568266 569894
rect 568502 569658 568586 569894
rect 568822 569658 568854 569894
rect 568234 569574 568854 569658
rect 568234 569338 568266 569574
rect 568502 569338 568586 569574
rect 568822 569338 568854 569574
rect 568234 533894 568854 569338
rect 568234 533658 568266 533894
rect 568502 533658 568586 533894
rect 568822 533658 568854 533894
rect 568234 533574 568854 533658
rect 568234 533338 568266 533574
rect 568502 533338 568586 533574
rect 568822 533338 568854 533574
rect 568234 497894 568854 533338
rect 568234 497658 568266 497894
rect 568502 497658 568586 497894
rect 568822 497658 568854 497894
rect 568234 497574 568854 497658
rect 568234 497338 568266 497574
rect 568502 497338 568586 497574
rect 568822 497338 568854 497574
rect 568234 461894 568854 497338
rect 568234 461658 568266 461894
rect 568502 461658 568586 461894
rect 568822 461658 568854 461894
rect 568234 461574 568854 461658
rect 568234 461338 568266 461574
rect 568502 461338 568586 461574
rect 568822 461338 568854 461574
rect 568234 425894 568854 461338
rect 568234 425658 568266 425894
rect 568502 425658 568586 425894
rect 568822 425658 568854 425894
rect 568234 425574 568854 425658
rect 568234 425338 568266 425574
rect 568502 425338 568586 425574
rect 568822 425338 568854 425574
rect 568234 389894 568854 425338
rect 568234 389658 568266 389894
rect 568502 389658 568586 389894
rect 568822 389658 568854 389894
rect 568234 389574 568854 389658
rect 568234 389338 568266 389574
rect 568502 389338 568586 389574
rect 568822 389338 568854 389574
rect 568234 353894 568854 389338
rect 568234 353658 568266 353894
rect 568502 353658 568586 353894
rect 568822 353658 568854 353894
rect 568234 353574 568854 353658
rect 568234 353338 568266 353574
rect 568502 353338 568586 353574
rect 568822 353338 568854 353574
rect 568234 317894 568854 353338
rect 568234 317658 568266 317894
rect 568502 317658 568586 317894
rect 568822 317658 568854 317894
rect 568234 317574 568854 317658
rect 568234 317338 568266 317574
rect 568502 317338 568586 317574
rect 568822 317338 568854 317574
rect 568234 281894 568854 317338
rect 568234 281658 568266 281894
rect 568502 281658 568586 281894
rect 568822 281658 568854 281894
rect 568234 281574 568854 281658
rect 568234 281338 568266 281574
rect 568502 281338 568586 281574
rect 568822 281338 568854 281574
rect 568234 245894 568854 281338
rect 568234 245658 568266 245894
rect 568502 245658 568586 245894
rect 568822 245658 568854 245894
rect 568234 245574 568854 245658
rect 568234 245338 568266 245574
rect 568502 245338 568586 245574
rect 568822 245338 568854 245574
rect 568234 209894 568854 245338
rect 568234 209658 568266 209894
rect 568502 209658 568586 209894
rect 568822 209658 568854 209894
rect 568234 209574 568854 209658
rect 568234 209338 568266 209574
rect 568502 209338 568586 209574
rect 568822 209338 568854 209574
rect 568234 173894 568854 209338
rect 568234 173658 568266 173894
rect 568502 173658 568586 173894
rect 568822 173658 568854 173894
rect 568234 173574 568854 173658
rect 568234 173338 568266 173574
rect 568502 173338 568586 173574
rect 568822 173338 568854 173574
rect 568234 137894 568854 173338
rect 568234 137658 568266 137894
rect 568502 137658 568586 137894
rect 568822 137658 568854 137894
rect 568234 137574 568854 137658
rect 568234 137338 568266 137574
rect 568502 137338 568586 137574
rect 568822 137338 568854 137574
rect 568234 101894 568854 137338
rect 568234 101658 568266 101894
rect 568502 101658 568586 101894
rect 568822 101658 568854 101894
rect 568234 101574 568854 101658
rect 568234 101338 568266 101574
rect 568502 101338 568586 101574
rect 568822 101338 568854 101574
rect 568234 65894 568854 101338
rect 568234 65658 568266 65894
rect 568502 65658 568586 65894
rect 568822 65658 568854 65894
rect 568234 65574 568854 65658
rect 568234 65338 568266 65574
rect 568502 65338 568586 65574
rect 568822 65338 568854 65574
rect 568234 29894 568854 65338
rect 568234 29658 568266 29894
rect 568502 29658 568586 29894
rect 568822 29658 568854 29894
rect 568234 29574 568854 29658
rect 568234 29338 568266 29574
rect 568502 29338 568586 29574
rect 568822 29338 568854 29574
rect 568234 -7066 568854 29338
rect 568234 -7302 568266 -7066
rect 568502 -7302 568586 -7066
rect 568822 -7302 568854 -7066
rect 568234 -7386 568854 -7302
rect 568234 -7622 568266 -7386
rect 568502 -7622 568586 -7386
rect 568822 -7622 568854 -7386
rect 568234 -7654 568854 -7622
rect 578194 704838 578814 711590
rect 578194 704602 578226 704838
rect 578462 704602 578546 704838
rect 578782 704602 578814 704838
rect 578194 704518 578814 704602
rect 578194 704282 578226 704518
rect 578462 704282 578546 704518
rect 578782 704282 578814 704518
rect 578194 687854 578814 704282
rect 578194 687618 578226 687854
rect 578462 687618 578546 687854
rect 578782 687618 578814 687854
rect 578194 687534 578814 687618
rect 578194 687298 578226 687534
rect 578462 687298 578546 687534
rect 578782 687298 578814 687534
rect 578194 651854 578814 687298
rect 578194 651618 578226 651854
rect 578462 651618 578546 651854
rect 578782 651618 578814 651854
rect 578194 651534 578814 651618
rect 578194 651298 578226 651534
rect 578462 651298 578546 651534
rect 578782 651298 578814 651534
rect 578194 615854 578814 651298
rect 578194 615618 578226 615854
rect 578462 615618 578546 615854
rect 578782 615618 578814 615854
rect 578194 615534 578814 615618
rect 578194 615298 578226 615534
rect 578462 615298 578546 615534
rect 578782 615298 578814 615534
rect 578194 579854 578814 615298
rect 578194 579618 578226 579854
rect 578462 579618 578546 579854
rect 578782 579618 578814 579854
rect 578194 579534 578814 579618
rect 578194 579298 578226 579534
rect 578462 579298 578546 579534
rect 578782 579298 578814 579534
rect 578194 543854 578814 579298
rect 578194 543618 578226 543854
rect 578462 543618 578546 543854
rect 578782 543618 578814 543854
rect 578194 543534 578814 543618
rect 578194 543298 578226 543534
rect 578462 543298 578546 543534
rect 578782 543298 578814 543534
rect 578194 507854 578814 543298
rect 578194 507618 578226 507854
rect 578462 507618 578546 507854
rect 578782 507618 578814 507854
rect 578194 507534 578814 507618
rect 578194 507298 578226 507534
rect 578462 507298 578546 507534
rect 578782 507298 578814 507534
rect 578194 471854 578814 507298
rect 578194 471618 578226 471854
rect 578462 471618 578546 471854
rect 578782 471618 578814 471854
rect 578194 471534 578814 471618
rect 578194 471298 578226 471534
rect 578462 471298 578546 471534
rect 578782 471298 578814 471534
rect 578194 435854 578814 471298
rect 578194 435618 578226 435854
rect 578462 435618 578546 435854
rect 578782 435618 578814 435854
rect 578194 435534 578814 435618
rect 578194 435298 578226 435534
rect 578462 435298 578546 435534
rect 578782 435298 578814 435534
rect 578194 399854 578814 435298
rect 578194 399618 578226 399854
rect 578462 399618 578546 399854
rect 578782 399618 578814 399854
rect 578194 399534 578814 399618
rect 578194 399298 578226 399534
rect 578462 399298 578546 399534
rect 578782 399298 578814 399534
rect 578194 363854 578814 399298
rect 578194 363618 578226 363854
rect 578462 363618 578546 363854
rect 578782 363618 578814 363854
rect 578194 363534 578814 363618
rect 578194 363298 578226 363534
rect 578462 363298 578546 363534
rect 578782 363298 578814 363534
rect 578194 327854 578814 363298
rect 578194 327618 578226 327854
rect 578462 327618 578546 327854
rect 578782 327618 578814 327854
rect 578194 327534 578814 327618
rect 578194 327298 578226 327534
rect 578462 327298 578546 327534
rect 578782 327298 578814 327534
rect 578194 291854 578814 327298
rect 578194 291618 578226 291854
rect 578462 291618 578546 291854
rect 578782 291618 578814 291854
rect 578194 291534 578814 291618
rect 578194 291298 578226 291534
rect 578462 291298 578546 291534
rect 578782 291298 578814 291534
rect 578194 255854 578814 291298
rect 578194 255618 578226 255854
rect 578462 255618 578546 255854
rect 578782 255618 578814 255854
rect 578194 255534 578814 255618
rect 578194 255298 578226 255534
rect 578462 255298 578546 255534
rect 578782 255298 578814 255534
rect 578194 219854 578814 255298
rect 578194 219618 578226 219854
rect 578462 219618 578546 219854
rect 578782 219618 578814 219854
rect 578194 219534 578814 219618
rect 578194 219298 578226 219534
rect 578462 219298 578546 219534
rect 578782 219298 578814 219534
rect 578194 183854 578814 219298
rect 578194 183618 578226 183854
rect 578462 183618 578546 183854
rect 578782 183618 578814 183854
rect 578194 183534 578814 183618
rect 578194 183298 578226 183534
rect 578462 183298 578546 183534
rect 578782 183298 578814 183534
rect 578194 147854 578814 183298
rect 578194 147618 578226 147854
rect 578462 147618 578546 147854
rect 578782 147618 578814 147854
rect 578194 147534 578814 147618
rect 578194 147298 578226 147534
rect 578462 147298 578546 147534
rect 578782 147298 578814 147534
rect 578194 111854 578814 147298
rect 578194 111618 578226 111854
rect 578462 111618 578546 111854
rect 578782 111618 578814 111854
rect 578194 111534 578814 111618
rect 578194 111298 578226 111534
rect 578462 111298 578546 111534
rect 578782 111298 578814 111534
rect 578194 75854 578814 111298
rect 578194 75618 578226 75854
rect 578462 75618 578546 75854
rect 578782 75618 578814 75854
rect 578194 75534 578814 75618
rect 578194 75298 578226 75534
rect 578462 75298 578546 75534
rect 578782 75298 578814 75534
rect 578194 39854 578814 75298
rect 578194 39618 578226 39854
rect 578462 39618 578546 39854
rect 578782 39618 578814 39854
rect 578194 39534 578814 39618
rect 578194 39298 578226 39534
rect 578462 39298 578546 39534
rect 578782 39298 578814 39534
rect 578194 3854 578814 39298
rect 578194 3618 578226 3854
rect 578462 3618 578546 3854
rect 578782 3618 578814 3854
rect 578194 3534 578814 3618
rect 578194 3298 578226 3534
rect 578462 3298 578546 3534
rect 578782 3298 578814 3534
rect 578194 -346 578814 3298
rect 578194 -582 578226 -346
rect 578462 -582 578546 -346
rect 578782 -582 578814 -346
rect 578194 -666 578814 -582
rect 578194 -902 578226 -666
rect 578462 -902 578546 -666
rect 578782 -902 578814 -666
rect 578194 -7654 578814 -902
rect 581914 705798 582534 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581914 705562 581946 705798
rect 582182 705562 582266 705798
rect 582502 705562 582534 705798
rect 581914 705478 582534 705562
rect 581914 705242 581946 705478
rect 582182 705242 582266 705478
rect 582502 705242 582534 705478
rect 581914 691574 582534 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581914 691338 581946 691574
rect 582182 691338 582266 691574
rect 582502 691338 582534 691574
rect 581914 691254 582534 691338
rect 581914 691018 581946 691254
rect 582182 691018 582266 691254
rect 582502 691018 582534 691254
rect 581914 655574 582534 691018
rect 581914 655338 581946 655574
rect 582182 655338 582266 655574
rect 582502 655338 582534 655574
rect 581914 655254 582534 655338
rect 581914 655018 581946 655254
rect 582182 655018 582266 655254
rect 582502 655018 582534 655254
rect 581914 619574 582534 655018
rect 581914 619338 581946 619574
rect 582182 619338 582266 619574
rect 582502 619338 582534 619574
rect 581914 619254 582534 619338
rect 581914 619018 581946 619254
rect 582182 619018 582266 619254
rect 582502 619018 582534 619254
rect 581914 583574 582534 619018
rect 581914 583338 581946 583574
rect 582182 583338 582266 583574
rect 582502 583338 582534 583574
rect 581914 583254 582534 583338
rect 581914 583018 581946 583254
rect 582182 583018 582266 583254
rect 582502 583018 582534 583254
rect 581914 547574 582534 583018
rect 581914 547338 581946 547574
rect 582182 547338 582266 547574
rect 582502 547338 582534 547574
rect 581914 547254 582534 547338
rect 581914 547018 581946 547254
rect 582182 547018 582266 547254
rect 582502 547018 582534 547254
rect 581914 511574 582534 547018
rect 581914 511338 581946 511574
rect 582182 511338 582266 511574
rect 582502 511338 582534 511574
rect 581914 511254 582534 511338
rect 581914 511018 581946 511254
rect 582182 511018 582266 511254
rect 582502 511018 582534 511254
rect 581914 475574 582534 511018
rect 581914 475338 581946 475574
rect 582182 475338 582266 475574
rect 582502 475338 582534 475574
rect 581914 475254 582534 475338
rect 581914 475018 581946 475254
rect 582182 475018 582266 475254
rect 582502 475018 582534 475254
rect 581914 439574 582534 475018
rect 581914 439338 581946 439574
rect 582182 439338 582266 439574
rect 582502 439338 582534 439574
rect 581914 439254 582534 439338
rect 581914 439018 581946 439254
rect 582182 439018 582266 439254
rect 582502 439018 582534 439254
rect 581914 403574 582534 439018
rect 581914 403338 581946 403574
rect 582182 403338 582266 403574
rect 582502 403338 582534 403574
rect 581914 403254 582534 403338
rect 581914 403018 581946 403254
rect 582182 403018 582266 403254
rect 582502 403018 582534 403254
rect 581914 367574 582534 403018
rect 581914 367338 581946 367574
rect 582182 367338 582266 367574
rect 582502 367338 582534 367574
rect 581914 367254 582534 367338
rect 581914 367018 581946 367254
rect 582182 367018 582266 367254
rect 582502 367018 582534 367254
rect 581914 331574 582534 367018
rect 581914 331338 581946 331574
rect 582182 331338 582266 331574
rect 582502 331338 582534 331574
rect 581914 331254 582534 331338
rect 581914 331018 581946 331254
rect 582182 331018 582266 331254
rect 582502 331018 582534 331254
rect 581914 295574 582534 331018
rect 581914 295338 581946 295574
rect 582182 295338 582266 295574
rect 582502 295338 582534 295574
rect 581914 295254 582534 295338
rect 581914 295018 581946 295254
rect 582182 295018 582266 295254
rect 582502 295018 582534 295254
rect 581914 259574 582534 295018
rect 581914 259338 581946 259574
rect 582182 259338 582266 259574
rect 582502 259338 582534 259574
rect 581914 259254 582534 259338
rect 581914 259018 581946 259254
rect 582182 259018 582266 259254
rect 582502 259018 582534 259254
rect 581914 223574 582534 259018
rect 581914 223338 581946 223574
rect 582182 223338 582266 223574
rect 582502 223338 582534 223574
rect 581914 223254 582534 223338
rect 581914 223018 581946 223254
rect 582182 223018 582266 223254
rect 582502 223018 582534 223254
rect 581914 187574 582534 223018
rect 581914 187338 581946 187574
rect 582182 187338 582266 187574
rect 582502 187338 582534 187574
rect 581914 187254 582534 187338
rect 581914 187018 581946 187254
rect 582182 187018 582266 187254
rect 582502 187018 582534 187254
rect 581914 151574 582534 187018
rect 581914 151338 581946 151574
rect 582182 151338 582266 151574
rect 582502 151338 582534 151574
rect 581914 151254 582534 151338
rect 581914 151018 581946 151254
rect 582182 151018 582266 151254
rect 582502 151018 582534 151254
rect 581914 115574 582534 151018
rect 581914 115338 581946 115574
rect 582182 115338 582266 115574
rect 582502 115338 582534 115574
rect 581914 115254 582534 115338
rect 581914 115018 581946 115254
rect 582182 115018 582266 115254
rect 582502 115018 582534 115254
rect 581914 79574 582534 115018
rect 581914 79338 581946 79574
rect 582182 79338 582266 79574
rect 582502 79338 582534 79574
rect 581914 79254 582534 79338
rect 581914 79018 581946 79254
rect 582182 79018 582266 79254
rect 582502 79018 582534 79254
rect 581914 43574 582534 79018
rect 581914 43338 581946 43574
rect 582182 43338 582266 43574
rect 582502 43338 582534 43574
rect 581914 43254 582534 43338
rect 581914 43018 581946 43254
rect 582182 43018 582266 43254
rect 582502 43018 582534 43254
rect 581914 7574 582534 43018
rect 581914 7338 581946 7574
rect 582182 7338 582266 7574
rect 582502 7338 582534 7574
rect 581914 7254 582534 7338
rect 581914 7018 581946 7254
rect 582182 7018 582266 7254
rect 582502 7018 582534 7254
rect 581914 -1306 582534 7018
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687854 585930 704282
rect 585310 687618 585342 687854
rect 585578 687618 585662 687854
rect 585898 687618 585930 687854
rect 585310 687534 585930 687618
rect 585310 687298 585342 687534
rect 585578 687298 585662 687534
rect 585898 687298 585930 687534
rect 585310 651854 585930 687298
rect 585310 651618 585342 651854
rect 585578 651618 585662 651854
rect 585898 651618 585930 651854
rect 585310 651534 585930 651618
rect 585310 651298 585342 651534
rect 585578 651298 585662 651534
rect 585898 651298 585930 651534
rect 585310 615854 585930 651298
rect 585310 615618 585342 615854
rect 585578 615618 585662 615854
rect 585898 615618 585930 615854
rect 585310 615534 585930 615618
rect 585310 615298 585342 615534
rect 585578 615298 585662 615534
rect 585898 615298 585930 615534
rect 585310 579854 585930 615298
rect 585310 579618 585342 579854
rect 585578 579618 585662 579854
rect 585898 579618 585930 579854
rect 585310 579534 585930 579618
rect 585310 579298 585342 579534
rect 585578 579298 585662 579534
rect 585898 579298 585930 579534
rect 585310 543854 585930 579298
rect 585310 543618 585342 543854
rect 585578 543618 585662 543854
rect 585898 543618 585930 543854
rect 585310 543534 585930 543618
rect 585310 543298 585342 543534
rect 585578 543298 585662 543534
rect 585898 543298 585930 543534
rect 585310 507854 585930 543298
rect 585310 507618 585342 507854
rect 585578 507618 585662 507854
rect 585898 507618 585930 507854
rect 585310 507534 585930 507618
rect 585310 507298 585342 507534
rect 585578 507298 585662 507534
rect 585898 507298 585930 507534
rect 585310 471854 585930 507298
rect 585310 471618 585342 471854
rect 585578 471618 585662 471854
rect 585898 471618 585930 471854
rect 585310 471534 585930 471618
rect 585310 471298 585342 471534
rect 585578 471298 585662 471534
rect 585898 471298 585930 471534
rect 585310 435854 585930 471298
rect 585310 435618 585342 435854
rect 585578 435618 585662 435854
rect 585898 435618 585930 435854
rect 585310 435534 585930 435618
rect 585310 435298 585342 435534
rect 585578 435298 585662 435534
rect 585898 435298 585930 435534
rect 585310 399854 585930 435298
rect 585310 399618 585342 399854
rect 585578 399618 585662 399854
rect 585898 399618 585930 399854
rect 585310 399534 585930 399618
rect 585310 399298 585342 399534
rect 585578 399298 585662 399534
rect 585898 399298 585930 399534
rect 585310 363854 585930 399298
rect 585310 363618 585342 363854
rect 585578 363618 585662 363854
rect 585898 363618 585930 363854
rect 585310 363534 585930 363618
rect 585310 363298 585342 363534
rect 585578 363298 585662 363534
rect 585898 363298 585930 363534
rect 585310 327854 585930 363298
rect 585310 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 585930 327854
rect 585310 327534 585930 327618
rect 585310 327298 585342 327534
rect 585578 327298 585662 327534
rect 585898 327298 585930 327534
rect 585310 291854 585930 327298
rect 585310 291618 585342 291854
rect 585578 291618 585662 291854
rect 585898 291618 585930 291854
rect 585310 291534 585930 291618
rect 585310 291298 585342 291534
rect 585578 291298 585662 291534
rect 585898 291298 585930 291534
rect 585310 255854 585930 291298
rect 585310 255618 585342 255854
rect 585578 255618 585662 255854
rect 585898 255618 585930 255854
rect 585310 255534 585930 255618
rect 585310 255298 585342 255534
rect 585578 255298 585662 255534
rect 585898 255298 585930 255534
rect 585310 219854 585930 255298
rect 585310 219618 585342 219854
rect 585578 219618 585662 219854
rect 585898 219618 585930 219854
rect 585310 219534 585930 219618
rect 585310 219298 585342 219534
rect 585578 219298 585662 219534
rect 585898 219298 585930 219534
rect 585310 183854 585930 219298
rect 585310 183618 585342 183854
rect 585578 183618 585662 183854
rect 585898 183618 585930 183854
rect 585310 183534 585930 183618
rect 585310 183298 585342 183534
rect 585578 183298 585662 183534
rect 585898 183298 585930 183534
rect 585310 147854 585930 183298
rect 585310 147618 585342 147854
rect 585578 147618 585662 147854
rect 585898 147618 585930 147854
rect 585310 147534 585930 147618
rect 585310 147298 585342 147534
rect 585578 147298 585662 147534
rect 585898 147298 585930 147534
rect 585310 111854 585930 147298
rect 585310 111618 585342 111854
rect 585578 111618 585662 111854
rect 585898 111618 585930 111854
rect 585310 111534 585930 111618
rect 585310 111298 585342 111534
rect 585578 111298 585662 111534
rect 585898 111298 585930 111534
rect 585310 75854 585930 111298
rect 585310 75618 585342 75854
rect 585578 75618 585662 75854
rect 585898 75618 585930 75854
rect 585310 75534 585930 75618
rect 585310 75298 585342 75534
rect 585578 75298 585662 75534
rect 585898 75298 585930 75534
rect 585310 39854 585930 75298
rect 585310 39618 585342 39854
rect 585578 39618 585662 39854
rect 585898 39618 585930 39854
rect 585310 39534 585930 39618
rect 585310 39298 585342 39534
rect 585578 39298 585662 39534
rect 585898 39298 585930 39534
rect 585310 3854 585930 39298
rect 585310 3618 585342 3854
rect 585578 3618 585662 3854
rect 585898 3618 585930 3854
rect 585310 3534 585930 3618
rect 585310 3298 585342 3534
rect 585578 3298 585662 3534
rect 585898 3298 585930 3534
rect 585310 -346 585930 3298
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691574 586890 705242
rect 586270 691338 586302 691574
rect 586538 691338 586622 691574
rect 586858 691338 586890 691574
rect 586270 691254 586890 691338
rect 586270 691018 586302 691254
rect 586538 691018 586622 691254
rect 586858 691018 586890 691254
rect 586270 655574 586890 691018
rect 586270 655338 586302 655574
rect 586538 655338 586622 655574
rect 586858 655338 586890 655574
rect 586270 655254 586890 655338
rect 586270 655018 586302 655254
rect 586538 655018 586622 655254
rect 586858 655018 586890 655254
rect 586270 619574 586890 655018
rect 586270 619338 586302 619574
rect 586538 619338 586622 619574
rect 586858 619338 586890 619574
rect 586270 619254 586890 619338
rect 586270 619018 586302 619254
rect 586538 619018 586622 619254
rect 586858 619018 586890 619254
rect 586270 583574 586890 619018
rect 586270 583338 586302 583574
rect 586538 583338 586622 583574
rect 586858 583338 586890 583574
rect 586270 583254 586890 583338
rect 586270 583018 586302 583254
rect 586538 583018 586622 583254
rect 586858 583018 586890 583254
rect 586270 547574 586890 583018
rect 586270 547338 586302 547574
rect 586538 547338 586622 547574
rect 586858 547338 586890 547574
rect 586270 547254 586890 547338
rect 586270 547018 586302 547254
rect 586538 547018 586622 547254
rect 586858 547018 586890 547254
rect 586270 511574 586890 547018
rect 586270 511338 586302 511574
rect 586538 511338 586622 511574
rect 586858 511338 586890 511574
rect 586270 511254 586890 511338
rect 586270 511018 586302 511254
rect 586538 511018 586622 511254
rect 586858 511018 586890 511254
rect 586270 475574 586890 511018
rect 586270 475338 586302 475574
rect 586538 475338 586622 475574
rect 586858 475338 586890 475574
rect 586270 475254 586890 475338
rect 586270 475018 586302 475254
rect 586538 475018 586622 475254
rect 586858 475018 586890 475254
rect 586270 439574 586890 475018
rect 586270 439338 586302 439574
rect 586538 439338 586622 439574
rect 586858 439338 586890 439574
rect 586270 439254 586890 439338
rect 586270 439018 586302 439254
rect 586538 439018 586622 439254
rect 586858 439018 586890 439254
rect 586270 403574 586890 439018
rect 586270 403338 586302 403574
rect 586538 403338 586622 403574
rect 586858 403338 586890 403574
rect 586270 403254 586890 403338
rect 586270 403018 586302 403254
rect 586538 403018 586622 403254
rect 586858 403018 586890 403254
rect 586270 367574 586890 403018
rect 586270 367338 586302 367574
rect 586538 367338 586622 367574
rect 586858 367338 586890 367574
rect 586270 367254 586890 367338
rect 586270 367018 586302 367254
rect 586538 367018 586622 367254
rect 586858 367018 586890 367254
rect 586270 331574 586890 367018
rect 586270 331338 586302 331574
rect 586538 331338 586622 331574
rect 586858 331338 586890 331574
rect 586270 331254 586890 331338
rect 586270 331018 586302 331254
rect 586538 331018 586622 331254
rect 586858 331018 586890 331254
rect 586270 295574 586890 331018
rect 586270 295338 586302 295574
rect 586538 295338 586622 295574
rect 586858 295338 586890 295574
rect 586270 295254 586890 295338
rect 586270 295018 586302 295254
rect 586538 295018 586622 295254
rect 586858 295018 586890 295254
rect 586270 259574 586890 295018
rect 586270 259338 586302 259574
rect 586538 259338 586622 259574
rect 586858 259338 586890 259574
rect 586270 259254 586890 259338
rect 586270 259018 586302 259254
rect 586538 259018 586622 259254
rect 586858 259018 586890 259254
rect 586270 223574 586890 259018
rect 586270 223338 586302 223574
rect 586538 223338 586622 223574
rect 586858 223338 586890 223574
rect 586270 223254 586890 223338
rect 586270 223018 586302 223254
rect 586538 223018 586622 223254
rect 586858 223018 586890 223254
rect 586270 187574 586890 223018
rect 586270 187338 586302 187574
rect 586538 187338 586622 187574
rect 586858 187338 586890 187574
rect 586270 187254 586890 187338
rect 586270 187018 586302 187254
rect 586538 187018 586622 187254
rect 586858 187018 586890 187254
rect 586270 151574 586890 187018
rect 586270 151338 586302 151574
rect 586538 151338 586622 151574
rect 586858 151338 586890 151574
rect 586270 151254 586890 151338
rect 586270 151018 586302 151254
rect 586538 151018 586622 151254
rect 586858 151018 586890 151254
rect 586270 115574 586890 151018
rect 586270 115338 586302 115574
rect 586538 115338 586622 115574
rect 586858 115338 586890 115574
rect 586270 115254 586890 115338
rect 586270 115018 586302 115254
rect 586538 115018 586622 115254
rect 586858 115018 586890 115254
rect 586270 79574 586890 115018
rect 586270 79338 586302 79574
rect 586538 79338 586622 79574
rect 586858 79338 586890 79574
rect 586270 79254 586890 79338
rect 586270 79018 586302 79254
rect 586538 79018 586622 79254
rect 586858 79018 586890 79254
rect 586270 43574 586890 79018
rect 586270 43338 586302 43574
rect 586538 43338 586622 43574
rect 586858 43338 586890 43574
rect 586270 43254 586890 43338
rect 586270 43018 586302 43254
rect 586538 43018 586622 43254
rect 586858 43018 586890 43254
rect 586270 7574 586890 43018
rect 586270 7338 586302 7574
rect 586538 7338 586622 7574
rect 586858 7338 586890 7574
rect 586270 7254 586890 7338
rect 586270 7018 586302 7254
rect 586538 7018 586622 7254
rect 586858 7018 586890 7254
rect 581914 -1542 581946 -1306
rect 582182 -1542 582266 -1306
rect 582502 -1542 582534 -1306
rect 581914 -1626 582534 -1542
rect 581914 -1862 581946 -1626
rect 582182 -1862 582266 -1626
rect 582502 -1862 582534 -1626
rect 581914 -7654 582534 -1862
rect 586270 -1306 586890 7018
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 695294 587850 706202
rect 587230 695058 587262 695294
rect 587498 695058 587582 695294
rect 587818 695058 587850 695294
rect 587230 694974 587850 695058
rect 587230 694738 587262 694974
rect 587498 694738 587582 694974
rect 587818 694738 587850 694974
rect 587230 659294 587850 694738
rect 587230 659058 587262 659294
rect 587498 659058 587582 659294
rect 587818 659058 587850 659294
rect 587230 658974 587850 659058
rect 587230 658738 587262 658974
rect 587498 658738 587582 658974
rect 587818 658738 587850 658974
rect 587230 623294 587850 658738
rect 587230 623058 587262 623294
rect 587498 623058 587582 623294
rect 587818 623058 587850 623294
rect 587230 622974 587850 623058
rect 587230 622738 587262 622974
rect 587498 622738 587582 622974
rect 587818 622738 587850 622974
rect 587230 587294 587850 622738
rect 587230 587058 587262 587294
rect 587498 587058 587582 587294
rect 587818 587058 587850 587294
rect 587230 586974 587850 587058
rect 587230 586738 587262 586974
rect 587498 586738 587582 586974
rect 587818 586738 587850 586974
rect 587230 551294 587850 586738
rect 587230 551058 587262 551294
rect 587498 551058 587582 551294
rect 587818 551058 587850 551294
rect 587230 550974 587850 551058
rect 587230 550738 587262 550974
rect 587498 550738 587582 550974
rect 587818 550738 587850 550974
rect 587230 515294 587850 550738
rect 587230 515058 587262 515294
rect 587498 515058 587582 515294
rect 587818 515058 587850 515294
rect 587230 514974 587850 515058
rect 587230 514738 587262 514974
rect 587498 514738 587582 514974
rect 587818 514738 587850 514974
rect 587230 479294 587850 514738
rect 587230 479058 587262 479294
rect 587498 479058 587582 479294
rect 587818 479058 587850 479294
rect 587230 478974 587850 479058
rect 587230 478738 587262 478974
rect 587498 478738 587582 478974
rect 587818 478738 587850 478974
rect 587230 443294 587850 478738
rect 587230 443058 587262 443294
rect 587498 443058 587582 443294
rect 587818 443058 587850 443294
rect 587230 442974 587850 443058
rect 587230 442738 587262 442974
rect 587498 442738 587582 442974
rect 587818 442738 587850 442974
rect 587230 407294 587850 442738
rect 587230 407058 587262 407294
rect 587498 407058 587582 407294
rect 587818 407058 587850 407294
rect 587230 406974 587850 407058
rect 587230 406738 587262 406974
rect 587498 406738 587582 406974
rect 587818 406738 587850 406974
rect 587230 371294 587850 406738
rect 587230 371058 587262 371294
rect 587498 371058 587582 371294
rect 587818 371058 587850 371294
rect 587230 370974 587850 371058
rect 587230 370738 587262 370974
rect 587498 370738 587582 370974
rect 587818 370738 587850 370974
rect 587230 335294 587850 370738
rect 587230 335058 587262 335294
rect 587498 335058 587582 335294
rect 587818 335058 587850 335294
rect 587230 334974 587850 335058
rect 587230 334738 587262 334974
rect 587498 334738 587582 334974
rect 587818 334738 587850 334974
rect 587230 299294 587850 334738
rect 587230 299058 587262 299294
rect 587498 299058 587582 299294
rect 587818 299058 587850 299294
rect 587230 298974 587850 299058
rect 587230 298738 587262 298974
rect 587498 298738 587582 298974
rect 587818 298738 587850 298974
rect 587230 263294 587850 298738
rect 587230 263058 587262 263294
rect 587498 263058 587582 263294
rect 587818 263058 587850 263294
rect 587230 262974 587850 263058
rect 587230 262738 587262 262974
rect 587498 262738 587582 262974
rect 587818 262738 587850 262974
rect 587230 227294 587850 262738
rect 587230 227058 587262 227294
rect 587498 227058 587582 227294
rect 587818 227058 587850 227294
rect 587230 226974 587850 227058
rect 587230 226738 587262 226974
rect 587498 226738 587582 226974
rect 587818 226738 587850 226974
rect 587230 191294 587850 226738
rect 587230 191058 587262 191294
rect 587498 191058 587582 191294
rect 587818 191058 587850 191294
rect 587230 190974 587850 191058
rect 587230 190738 587262 190974
rect 587498 190738 587582 190974
rect 587818 190738 587850 190974
rect 587230 155294 587850 190738
rect 587230 155058 587262 155294
rect 587498 155058 587582 155294
rect 587818 155058 587850 155294
rect 587230 154974 587850 155058
rect 587230 154738 587262 154974
rect 587498 154738 587582 154974
rect 587818 154738 587850 154974
rect 587230 119294 587850 154738
rect 587230 119058 587262 119294
rect 587498 119058 587582 119294
rect 587818 119058 587850 119294
rect 587230 118974 587850 119058
rect 587230 118738 587262 118974
rect 587498 118738 587582 118974
rect 587818 118738 587850 118974
rect 587230 83294 587850 118738
rect 587230 83058 587262 83294
rect 587498 83058 587582 83294
rect 587818 83058 587850 83294
rect 587230 82974 587850 83058
rect 587230 82738 587262 82974
rect 587498 82738 587582 82974
rect 587818 82738 587850 82974
rect 587230 47294 587850 82738
rect 587230 47058 587262 47294
rect 587498 47058 587582 47294
rect 587818 47058 587850 47294
rect 587230 46974 587850 47058
rect 587230 46738 587262 46974
rect 587498 46738 587582 46974
rect 587818 46738 587850 46974
rect 587230 11294 587850 46738
rect 587230 11058 587262 11294
rect 587498 11058 587582 11294
rect 587818 11058 587850 11294
rect 587230 10974 587850 11058
rect 587230 10738 587262 10974
rect 587498 10738 587582 10974
rect 587818 10738 587850 10974
rect 587230 -2266 587850 10738
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 699014 588810 707162
rect 588190 698778 588222 699014
rect 588458 698778 588542 699014
rect 588778 698778 588810 699014
rect 588190 698694 588810 698778
rect 588190 698458 588222 698694
rect 588458 698458 588542 698694
rect 588778 698458 588810 698694
rect 588190 663014 588810 698458
rect 588190 662778 588222 663014
rect 588458 662778 588542 663014
rect 588778 662778 588810 663014
rect 588190 662694 588810 662778
rect 588190 662458 588222 662694
rect 588458 662458 588542 662694
rect 588778 662458 588810 662694
rect 588190 627014 588810 662458
rect 588190 626778 588222 627014
rect 588458 626778 588542 627014
rect 588778 626778 588810 627014
rect 588190 626694 588810 626778
rect 588190 626458 588222 626694
rect 588458 626458 588542 626694
rect 588778 626458 588810 626694
rect 588190 591014 588810 626458
rect 588190 590778 588222 591014
rect 588458 590778 588542 591014
rect 588778 590778 588810 591014
rect 588190 590694 588810 590778
rect 588190 590458 588222 590694
rect 588458 590458 588542 590694
rect 588778 590458 588810 590694
rect 588190 555014 588810 590458
rect 588190 554778 588222 555014
rect 588458 554778 588542 555014
rect 588778 554778 588810 555014
rect 588190 554694 588810 554778
rect 588190 554458 588222 554694
rect 588458 554458 588542 554694
rect 588778 554458 588810 554694
rect 588190 519014 588810 554458
rect 588190 518778 588222 519014
rect 588458 518778 588542 519014
rect 588778 518778 588810 519014
rect 588190 518694 588810 518778
rect 588190 518458 588222 518694
rect 588458 518458 588542 518694
rect 588778 518458 588810 518694
rect 588190 483014 588810 518458
rect 588190 482778 588222 483014
rect 588458 482778 588542 483014
rect 588778 482778 588810 483014
rect 588190 482694 588810 482778
rect 588190 482458 588222 482694
rect 588458 482458 588542 482694
rect 588778 482458 588810 482694
rect 588190 447014 588810 482458
rect 588190 446778 588222 447014
rect 588458 446778 588542 447014
rect 588778 446778 588810 447014
rect 588190 446694 588810 446778
rect 588190 446458 588222 446694
rect 588458 446458 588542 446694
rect 588778 446458 588810 446694
rect 588190 411014 588810 446458
rect 588190 410778 588222 411014
rect 588458 410778 588542 411014
rect 588778 410778 588810 411014
rect 588190 410694 588810 410778
rect 588190 410458 588222 410694
rect 588458 410458 588542 410694
rect 588778 410458 588810 410694
rect 588190 375014 588810 410458
rect 588190 374778 588222 375014
rect 588458 374778 588542 375014
rect 588778 374778 588810 375014
rect 588190 374694 588810 374778
rect 588190 374458 588222 374694
rect 588458 374458 588542 374694
rect 588778 374458 588810 374694
rect 588190 339014 588810 374458
rect 588190 338778 588222 339014
rect 588458 338778 588542 339014
rect 588778 338778 588810 339014
rect 588190 338694 588810 338778
rect 588190 338458 588222 338694
rect 588458 338458 588542 338694
rect 588778 338458 588810 338694
rect 588190 303014 588810 338458
rect 588190 302778 588222 303014
rect 588458 302778 588542 303014
rect 588778 302778 588810 303014
rect 588190 302694 588810 302778
rect 588190 302458 588222 302694
rect 588458 302458 588542 302694
rect 588778 302458 588810 302694
rect 588190 267014 588810 302458
rect 588190 266778 588222 267014
rect 588458 266778 588542 267014
rect 588778 266778 588810 267014
rect 588190 266694 588810 266778
rect 588190 266458 588222 266694
rect 588458 266458 588542 266694
rect 588778 266458 588810 266694
rect 588190 231014 588810 266458
rect 588190 230778 588222 231014
rect 588458 230778 588542 231014
rect 588778 230778 588810 231014
rect 588190 230694 588810 230778
rect 588190 230458 588222 230694
rect 588458 230458 588542 230694
rect 588778 230458 588810 230694
rect 588190 195014 588810 230458
rect 588190 194778 588222 195014
rect 588458 194778 588542 195014
rect 588778 194778 588810 195014
rect 588190 194694 588810 194778
rect 588190 194458 588222 194694
rect 588458 194458 588542 194694
rect 588778 194458 588810 194694
rect 588190 159014 588810 194458
rect 588190 158778 588222 159014
rect 588458 158778 588542 159014
rect 588778 158778 588810 159014
rect 588190 158694 588810 158778
rect 588190 158458 588222 158694
rect 588458 158458 588542 158694
rect 588778 158458 588810 158694
rect 588190 123014 588810 158458
rect 588190 122778 588222 123014
rect 588458 122778 588542 123014
rect 588778 122778 588810 123014
rect 588190 122694 588810 122778
rect 588190 122458 588222 122694
rect 588458 122458 588542 122694
rect 588778 122458 588810 122694
rect 588190 87014 588810 122458
rect 588190 86778 588222 87014
rect 588458 86778 588542 87014
rect 588778 86778 588810 87014
rect 588190 86694 588810 86778
rect 588190 86458 588222 86694
rect 588458 86458 588542 86694
rect 588778 86458 588810 86694
rect 588190 51014 588810 86458
rect 588190 50778 588222 51014
rect 588458 50778 588542 51014
rect 588778 50778 588810 51014
rect 588190 50694 588810 50778
rect 588190 50458 588222 50694
rect 588458 50458 588542 50694
rect 588778 50458 588810 50694
rect 588190 15014 588810 50458
rect 588190 14778 588222 15014
rect 588458 14778 588542 15014
rect 588778 14778 588810 15014
rect 588190 14694 588810 14778
rect 588190 14458 588222 14694
rect 588458 14458 588542 14694
rect 588778 14458 588810 14694
rect 588190 -3226 588810 14458
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666734 589770 708122
rect 589150 666498 589182 666734
rect 589418 666498 589502 666734
rect 589738 666498 589770 666734
rect 589150 666414 589770 666498
rect 589150 666178 589182 666414
rect 589418 666178 589502 666414
rect 589738 666178 589770 666414
rect 589150 630734 589770 666178
rect 589150 630498 589182 630734
rect 589418 630498 589502 630734
rect 589738 630498 589770 630734
rect 589150 630414 589770 630498
rect 589150 630178 589182 630414
rect 589418 630178 589502 630414
rect 589738 630178 589770 630414
rect 589150 594734 589770 630178
rect 589150 594498 589182 594734
rect 589418 594498 589502 594734
rect 589738 594498 589770 594734
rect 589150 594414 589770 594498
rect 589150 594178 589182 594414
rect 589418 594178 589502 594414
rect 589738 594178 589770 594414
rect 589150 558734 589770 594178
rect 589150 558498 589182 558734
rect 589418 558498 589502 558734
rect 589738 558498 589770 558734
rect 589150 558414 589770 558498
rect 589150 558178 589182 558414
rect 589418 558178 589502 558414
rect 589738 558178 589770 558414
rect 589150 522734 589770 558178
rect 589150 522498 589182 522734
rect 589418 522498 589502 522734
rect 589738 522498 589770 522734
rect 589150 522414 589770 522498
rect 589150 522178 589182 522414
rect 589418 522178 589502 522414
rect 589738 522178 589770 522414
rect 589150 486734 589770 522178
rect 589150 486498 589182 486734
rect 589418 486498 589502 486734
rect 589738 486498 589770 486734
rect 589150 486414 589770 486498
rect 589150 486178 589182 486414
rect 589418 486178 589502 486414
rect 589738 486178 589770 486414
rect 589150 450734 589770 486178
rect 589150 450498 589182 450734
rect 589418 450498 589502 450734
rect 589738 450498 589770 450734
rect 589150 450414 589770 450498
rect 589150 450178 589182 450414
rect 589418 450178 589502 450414
rect 589738 450178 589770 450414
rect 589150 414734 589770 450178
rect 589150 414498 589182 414734
rect 589418 414498 589502 414734
rect 589738 414498 589770 414734
rect 589150 414414 589770 414498
rect 589150 414178 589182 414414
rect 589418 414178 589502 414414
rect 589738 414178 589770 414414
rect 589150 378734 589770 414178
rect 589150 378498 589182 378734
rect 589418 378498 589502 378734
rect 589738 378498 589770 378734
rect 589150 378414 589770 378498
rect 589150 378178 589182 378414
rect 589418 378178 589502 378414
rect 589738 378178 589770 378414
rect 589150 342734 589770 378178
rect 589150 342498 589182 342734
rect 589418 342498 589502 342734
rect 589738 342498 589770 342734
rect 589150 342414 589770 342498
rect 589150 342178 589182 342414
rect 589418 342178 589502 342414
rect 589738 342178 589770 342414
rect 589150 306734 589770 342178
rect 589150 306498 589182 306734
rect 589418 306498 589502 306734
rect 589738 306498 589770 306734
rect 589150 306414 589770 306498
rect 589150 306178 589182 306414
rect 589418 306178 589502 306414
rect 589738 306178 589770 306414
rect 589150 270734 589770 306178
rect 589150 270498 589182 270734
rect 589418 270498 589502 270734
rect 589738 270498 589770 270734
rect 589150 270414 589770 270498
rect 589150 270178 589182 270414
rect 589418 270178 589502 270414
rect 589738 270178 589770 270414
rect 589150 234734 589770 270178
rect 589150 234498 589182 234734
rect 589418 234498 589502 234734
rect 589738 234498 589770 234734
rect 589150 234414 589770 234498
rect 589150 234178 589182 234414
rect 589418 234178 589502 234414
rect 589738 234178 589770 234414
rect 589150 198734 589770 234178
rect 589150 198498 589182 198734
rect 589418 198498 589502 198734
rect 589738 198498 589770 198734
rect 589150 198414 589770 198498
rect 589150 198178 589182 198414
rect 589418 198178 589502 198414
rect 589738 198178 589770 198414
rect 589150 162734 589770 198178
rect 589150 162498 589182 162734
rect 589418 162498 589502 162734
rect 589738 162498 589770 162734
rect 589150 162414 589770 162498
rect 589150 162178 589182 162414
rect 589418 162178 589502 162414
rect 589738 162178 589770 162414
rect 589150 126734 589770 162178
rect 589150 126498 589182 126734
rect 589418 126498 589502 126734
rect 589738 126498 589770 126734
rect 589150 126414 589770 126498
rect 589150 126178 589182 126414
rect 589418 126178 589502 126414
rect 589738 126178 589770 126414
rect 589150 90734 589770 126178
rect 589150 90498 589182 90734
rect 589418 90498 589502 90734
rect 589738 90498 589770 90734
rect 589150 90414 589770 90498
rect 589150 90178 589182 90414
rect 589418 90178 589502 90414
rect 589738 90178 589770 90414
rect 589150 54734 589770 90178
rect 589150 54498 589182 54734
rect 589418 54498 589502 54734
rect 589738 54498 589770 54734
rect 589150 54414 589770 54498
rect 589150 54178 589182 54414
rect 589418 54178 589502 54414
rect 589738 54178 589770 54414
rect 589150 18734 589770 54178
rect 589150 18498 589182 18734
rect 589418 18498 589502 18734
rect 589738 18498 589770 18734
rect 589150 18414 589770 18498
rect 589150 18178 589182 18414
rect 589418 18178 589502 18414
rect 589738 18178 589770 18414
rect 589150 -4186 589770 18178
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670454 590730 709082
rect 590110 670218 590142 670454
rect 590378 670218 590462 670454
rect 590698 670218 590730 670454
rect 590110 670134 590730 670218
rect 590110 669898 590142 670134
rect 590378 669898 590462 670134
rect 590698 669898 590730 670134
rect 590110 634454 590730 669898
rect 590110 634218 590142 634454
rect 590378 634218 590462 634454
rect 590698 634218 590730 634454
rect 590110 634134 590730 634218
rect 590110 633898 590142 634134
rect 590378 633898 590462 634134
rect 590698 633898 590730 634134
rect 590110 598454 590730 633898
rect 590110 598218 590142 598454
rect 590378 598218 590462 598454
rect 590698 598218 590730 598454
rect 590110 598134 590730 598218
rect 590110 597898 590142 598134
rect 590378 597898 590462 598134
rect 590698 597898 590730 598134
rect 590110 562454 590730 597898
rect 590110 562218 590142 562454
rect 590378 562218 590462 562454
rect 590698 562218 590730 562454
rect 590110 562134 590730 562218
rect 590110 561898 590142 562134
rect 590378 561898 590462 562134
rect 590698 561898 590730 562134
rect 590110 526454 590730 561898
rect 590110 526218 590142 526454
rect 590378 526218 590462 526454
rect 590698 526218 590730 526454
rect 590110 526134 590730 526218
rect 590110 525898 590142 526134
rect 590378 525898 590462 526134
rect 590698 525898 590730 526134
rect 590110 490454 590730 525898
rect 590110 490218 590142 490454
rect 590378 490218 590462 490454
rect 590698 490218 590730 490454
rect 590110 490134 590730 490218
rect 590110 489898 590142 490134
rect 590378 489898 590462 490134
rect 590698 489898 590730 490134
rect 590110 454454 590730 489898
rect 590110 454218 590142 454454
rect 590378 454218 590462 454454
rect 590698 454218 590730 454454
rect 590110 454134 590730 454218
rect 590110 453898 590142 454134
rect 590378 453898 590462 454134
rect 590698 453898 590730 454134
rect 590110 418454 590730 453898
rect 590110 418218 590142 418454
rect 590378 418218 590462 418454
rect 590698 418218 590730 418454
rect 590110 418134 590730 418218
rect 590110 417898 590142 418134
rect 590378 417898 590462 418134
rect 590698 417898 590730 418134
rect 590110 382454 590730 417898
rect 590110 382218 590142 382454
rect 590378 382218 590462 382454
rect 590698 382218 590730 382454
rect 590110 382134 590730 382218
rect 590110 381898 590142 382134
rect 590378 381898 590462 382134
rect 590698 381898 590730 382134
rect 590110 346454 590730 381898
rect 590110 346218 590142 346454
rect 590378 346218 590462 346454
rect 590698 346218 590730 346454
rect 590110 346134 590730 346218
rect 590110 345898 590142 346134
rect 590378 345898 590462 346134
rect 590698 345898 590730 346134
rect 590110 310454 590730 345898
rect 590110 310218 590142 310454
rect 590378 310218 590462 310454
rect 590698 310218 590730 310454
rect 590110 310134 590730 310218
rect 590110 309898 590142 310134
rect 590378 309898 590462 310134
rect 590698 309898 590730 310134
rect 590110 274454 590730 309898
rect 590110 274218 590142 274454
rect 590378 274218 590462 274454
rect 590698 274218 590730 274454
rect 590110 274134 590730 274218
rect 590110 273898 590142 274134
rect 590378 273898 590462 274134
rect 590698 273898 590730 274134
rect 590110 238454 590730 273898
rect 590110 238218 590142 238454
rect 590378 238218 590462 238454
rect 590698 238218 590730 238454
rect 590110 238134 590730 238218
rect 590110 237898 590142 238134
rect 590378 237898 590462 238134
rect 590698 237898 590730 238134
rect 590110 202454 590730 237898
rect 590110 202218 590142 202454
rect 590378 202218 590462 202454
rect 590698 202218 590730 202454
rect 590110 202134 590730 202218
rect 590110 201898 590142 202134
rect 590378 201898 590462 202134
rect 590698 201898 590730 202134
rect 590110 166454 590730 201898
rect 590110 166218 590142 166454
rect 590378 166218 590462 166454
rect 590698 166218 590730 166454
rect 590110 166134 590730 166218
rect 590110 165898 590142 166134
rect 590378 165898 590462 166134
rect 590698 165898 590730 166134
rect 590110 130454 590730 165898
rect 590110 130218 590142 130454
rect 590378 130218 590462 130454
rect 590698 130218 590730 130454
rect 590110 130134 590730 130218
rect 590110 129898 590142 130134
rect 590378 129898 590462 130134
rect 590698 129898 590730 130134
rect 590110 94454 590730 129898
rect 590110 94218 590142 94454
rect 590378 94218 590462 94454
rect 590698 94218 590730 94454
rect 590110 94134 590730 94218
rect 590110 93898 590142 94134
rect 590378 93898 590462 94134
rect 590698 93898 590730 94134
rect 590110 58454 590730 93898
rect 590110 58218 590142 58454
rect 590378 58218 590462 58454
rect 590698 58218 590730 58454
rect 590110 58134 590730 58218
rect 590110 57898 590142 58134
rect 590378 57898 590462 58134
rect 590698 57898 590730 58134
rect 590110 22454 590730 57898
rect 590110 22218 590142 22454
rect 590378 22218 590462 22454
rect 590698 22218 590730 22454
rect 590110 22134 590730 22218
rect 590110 21898 590142 22134
rect 590378 21898 590462 22134
rect 590698 21898 590730 22134
rect 590110 -5146 590730 21898
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 674174 591690 710042
rect 591070 673938 591102 674174
rect 591338 673938 591422 674174
rect 591658 673938 591690 674174
rect 591070 673854 591690 673938
rect 591070 673618 591102 673854
rect 591338 673618 591422 673854
rect 591658 673618 591690 673854
rect 591070 638174 591690 673618
rect 591070 637938 591102 638174
rect 591338 637938 591422 638174
rect 591658 637938 591690 638174
rect 591070 637854 591690 637938
rect 591070 637618 591102 637854
rect 591338 637618 591422 637854
rect 591658 637618 591690 637854
rect 591070 602174 591690 637618
rect 591070 601938 591102 602174
rect 591338 601938 591422 602174
rect 591658 601938 591690 602174
rect 591070 601854 591690 601938
rect 591070 601618 591102 601854
rect 591338 601618 591422 601854
rect 591658 601618 591690 601854
rect 591070 566174 591690 601618
rect 591070 565938 591102 566174
rect 591338 565938 591422 566174
rect 591658 565938 591690 566174
rect 591070 565854 591690 565938
rect 591070 565618 591102 565854
rect 591338 565618 591422 565854
rect 591658 565618 591690 565854
rect 591070 530174 591690 565618
rect 591070 529938 591102 530174
rect 591338 529938 591422 530174
rect 591658 529938 591690 530174
rect 591070 529854 591690 529938
rect 591070 529618 591102 529854
rect 591338 529618 591422 529854
rect 591658 529618 591690 529854
rect 591070 494174 591690 529618
rect 591070 493938 591102 494174
rect 591338 493938 591422 494174
rect 591658 493938 591690 494174
rect 591070 493854 591690 493938
rect 591070 493618 591102 493854
rect 591338 493618 591422 493854
rect 591658 493618 591690 493854
rect 591070 458174 591690 493618
rect 591070 457938 591102 458174
rect 591338 457938 591422 458174
rect 591658 457938 591690 458174
rect 591070 457854 591690 457938
rect 591070 457618 591102 457854
rect 591338 457618 591422 457854
rect 591658 457618 591690 457854
rect 591070 422174 591690 457618
rect 591070 421938 591102 422174
rect 591338 421938 591422 422174
rect 591658 421938 591690 422174
rect 591070 421854 591690 421938
rect 591070 421618 591102 421854
rect 591338 421618 591422 421854
rect 591658 421618 591690 421854
rect 591070 386174 591690 421618
rect 591070 385938 591102 386174
rect 591338 385938 591422 386174
rect 591658 385938 591690 386174
rect 591070 385854 591690 385938
rect 591070 385618 591102 385854
rect 591338 385618 591422 385854
rect 591658 385618 591690 385854
rect 591070 350174 591690 385618
rect 591070 349938 591102 350174
rect 591338 349938 591422 350174
rect 591658 349938 591690 350174
rect 591070 349854 591690 349938
rect 591070 349618 591102 349854
rect 591338 349618 591422 349854
rect 591658 349618 591690 349854
rect 591070 314174 591690 349618
rect 591070 313938 591102 314174
rect 591338 313938 591422 314174
rect 591658 313938 591690 314174
rect 591070 313854 591690 313938
rect 591070 313618 591102 313854
rect 591338 313618 591422 313854
rect 591658 313618 591690 313854
rect 591070 278174 591690 313618
rect 591070 277938 591102 278174
rect 591338 277938 591422 278174
rect 591658 277938 591690 278174
rect 591070 277854 591690 277938
rect 591070 277618 591102 277854
rect 591338 277618 591422 277854
rect 591658 277618 591690 277854
rect 591070 242174 591690 277618
rect 591070 241938 591102 242174
rect 591338 241938 591422 242174
rect 591658 241938 591690 242174
rect 591070 241854 591690 241938
rect 591070 241618 591102 241854
rect 591338 241618 591422 241854
rect 591658 241618 591690 241854
rect 591070 206174 591690 241618
rect 591070 205938 591102 206174
rect 591338 205938 591422 206174
rect 591658 205938 591690 206174
rect 591070 205854 591690 205938
rect 591070 205618 591102 205854
rect 591338 205618 591422 205854
rect 591658 205618 591690 205854
rect 591070 170174 591690 205618
rect 591070 169938 591102 170174
rect 591338 169938 591422 170174
rect 591658 169938 591690 170174
rect 591070 169854 591690 169938
rect 591070 169618 591102 169854
rect 591338 169618 591422 169854
rect 591658 169618 591690 169854
rect 591070 134174 591690 169618
rect 591070 133938 591102 134174
rect 591338 133938 591422 134174
rect 591658 133938 591690 134174
rect 591070 133854 591690 133938
rect 591070 133618 591102 133854
rect 591338 133618 591422 133854
rect 591658 133618 591690 133854
rect 591070 98174 591690 133618
rect 591070 97938 591102 98174
rect 591338 97938 591422 98174
rect 591658 97938 591690 98174
rect 591070 97854 591690 97938
rect 591070 97618 591102 97854
rect 591338 97618 591422 97854
rect 591658 97618 591690 97854
rect 591070 62174 591690 97618
rect 591070 61938 591102 62174
rect 591338 61938 591422 62174
rect 591658 61938 591690 62174
rect 591070 61854 591690 61938
rect 591070 61618 591102 61854
rect 591338 61618 591422 61854
rect 591658 61618 591690 61854
rect 591070 26174 591690 61618
rect 591070 25938 591102 26174
rect 591338 25938 591422 26174
rect 591658 25938 591690 26174
rect 591070 25854 591690 25938
rect 591070 25618 591102 25854
rect 591338 25618 591422 25854
rect 591658 25618 591690 25854
rect 591070 -6106 591690 25618
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677894 592650 711002
rect 592030 677658 592062 677894
rect 592298 677658 592382 677894
rect 592618 677658 592650 677894
rect 592030 677574 592650 677658
rect 592030 677338 592062 677574
rect 592298 677338 592382 677574
rect 592618 677338 592650 677574
rect 592030 641894 592650 677338
rect 592030 641658 592062 641894
rect 592298 641658 592382 641894
rect 592618 641658 592650 641894
rect 592030 641574 592650 641658
rect 592030 641338 592062 641574
rect 592298 641338 592382 641574
rect 592618 641338 592650 641574
rect 592030 605894 592650 641338
rect 592030 605658 592062 605894
rect 592298 605658 592382 605894
rect 592618 605658 592650 605894
rect 592030 605574 592650 605658
rect 592030 605338 592062 605574
rect 592298 605338 592382 605574
rect 592618 605338 592650 605574
rect 592030 569894 592650 605338
rect 592030 569658 592062 569894
rect 592298 569658 592382 569894
rect 592618 569658 592650 569894
rect 592030 569574 592650 569658
rect 592030 569338 592062 569574
rect 592298 569338 592382 569574
rect 592618 569338 592650 569574
rect 592030 533894 592650 569338
rect 592030 533658 592062 533894
rect 592298 533658 592382 533894
rect 592618 533658 592650 533894
rect 592030 533574 592650 533658
rect 592030 533338 592062 533574
rect 592298 533338 592382 533574
rect 592618 533338 592650 533574
rect 592030 497894 592650 533338
rect 592030 497658 592062 497894
rect 592298 497658 592382 497894
rect 592618 497658 592650 497894
rect 592030 497574 592650 497658
rect 592030 497338 592062 497574
rect 592298 497338 592382 497574
rect 592618 497338 592650 497574
rect 592030 461894 592650 497338
rect 592030 461658 592062 461894
rect 592298 461658 592382 461894
rect 592618 461658 592650 461894
rect 592030 461574 592650 461658
rect 592030 461338 592062 461574
rect 592298 461338 592382 461574
rect 592618 461338 592650 461574
rect 592030 425894 592650 461338
rect 592030 425658 592062 425894
rect 592298 425658 592382 425894
rect 592618 425658 592650 425894
rect 592030 425574 592650 425658
rect 592030 425338 592062 425574
rect 592298 425338 592382 425574
rect 592618 425338 592650 425574
rect 592030 389894 592650 425338
rect 592030 389658 592062 389894
rect 592298 389658 592382 389894
rect 592618 389658 592650 389894
rect 592030 389574 592650 389658
rect 592030 389338 592062 389574
rect 592298 389338 592382 389574
rect 592618 389338 592650 389574
rect 592030 353894 592650 389338
rect 592030 353658 592062 353894
rect 592298 353658 592382 353894
rect 592618 353658 592650 353894
rect 592030 353574 592650 353658
rect 592030 353338 592062 353574
rect 592298 353338 592382 353574
rect 592618 353338 592650 353574
rect 592030 317894 592650 353338
rect 592030 317658 592062 317894
rect 592298 317658 592382 317894
rect 592618 317658 592650 317894
rect 592030 317574 592650 317658
rect 592030 317338 592062 317574
rect 592298 317338 592382 317574
rect 592618 317338 592650 317574
rect 592030 281894 592650 317338
rect 592030 281658 592062 281894
rect 592298 281658 592382 281894
rect 592618 281658 592650 281894
rect 592030 281574 592650 281658
rect 592030 281338 592062 281574
rect 592298 281338 592382 281574
rect 592618 281338 592650 281574
rect 592030 245894 592650 281338
rect 592030 245658 592062 245894
rect 592298 245658 592382 245894
rect 592618 245658 592650 245894
rect 592030 245574 592650 245658
rect 592030 245338 592062 245574
rect 592298 245338 592382 245574
rect 592618 245338 592650 245574
rect 592030 209894 592650 245338
rect 592030 209658 592062 209894
rect 592298 209658 592382 209894
rect 592618 209658 592650 209894
rect 592030 209574 592650 209658
rect 592030 209338 592062 209574
rect 592298 209338 592382 209574
rect 592618 209338 592650 209574
rect 592030 173894 592650 209338
rect 592030 173658 592062 173894
rect 592298 173658 592382 173894
rect 592618 173658 592650 173894
rect 592030 173574 592650 173658
rect 592030 173338 592062 173574
rect 592298 173338 592382 173574
rect 592618 173338 592650 173574
rect 592030 137894 592650 173338
rect 592030 137658 592062 137894
rect 592298 137658 592382 137894
rect 592618 137658 592650 137894
rect 592030 137574 592650 137658
rect 592030 137338 592062 137574
rect 592298 137338 592382 137574
rect 592618 137338 592650 137574
rect 592030 101894 592650 137338
rect 592030 101658 592062 101894
rect 592298 101658 592382 101894
rect 592618 101658 592650 101894
rect 592030 101574 592650 101658
rect 592030 101338 592062 101574
rect 592298 101338 592382 101574
rect 592618 101338 592650 101574
rect 592030 65894 592650 101338
rect 592030 65658 592062 65894
rect 592298 65658 592382 65894
rect 592618 65658 592650 65894
rect 592030 65574 592650 65658
rect 592030 65338 592062 65574
rect 592298 65338 592382 65574
rect 592618 65338 592650 65574
rect 592030 29894 592650 65338
rect 592030 29658 592062 29894
rect 592298 29658 592382 29894
rect 592618 29658 592650 29894
rect 592030 29574 592650 29658
rect 592030 29338 592062 29574
rect 592298 29338 592382 29574
rect 592618 29338 592650 29574
rect 592030 -7066 592650 29338
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677658 -8458 677894
rect -8374 677658 -8138 677894
rect -8694 677338 -8458 677574
rect -8374 677338 -8138 677574
rect -8694 641658 -8458 641894
rect -8374 641658 -8138 641894
rect -8694 641338 -8458 641574
rect -8374 641338 -8138 641574
rect -8694 605658 -8458 605894
rect -8374 605658 -8138 605894
rect -8694 605338 -8458 605574
rect -8374 605338 -8138 605574
rect -8694 569658 -8458 569894
rect -8374 569658 -8138 569894
rect -8694 569338 -8458 569574
rect -8374 569338 -8138 569574
rect -8694 533658 -8458 533894
rect -8374 533658 -8138 533894
rect -8694 533338 -8458 533574
rect -8374 533338 -8138 533574
rect -8694 497658 -8458 497894
rect -8374 497658 -8138 497894
rect -8694 497338 -8458 497574
rect -8374 497338 -8138 497574
rect -8694 461658 -8458 461894
rect -8374 461658 -8138 461894
rect -8694 461338 -8458 461574
rect -8374 461338 -8138 461574
rect -8694 425658 -8458 425894
rect -8374 425658 -8138 425894
rect -8694 425338 -8458 425574
rect -8374 425338 -8138 425574
rect -8694 389658 -8458 389894
rect -8374 389658 -8138 389894
rect -8694 389338 -8458 389574
rect -8374 389338 -8138 389574
rect -8694 353658 -8458 353894
rect -8374 353658 -8138 353894
rect -8694 353338 -8458 353574
rect -8374 353338 -8138 353574
rect -8694 317658 -8458 317894
rect -8374 317658 -8138 317894
rect -8694 317338 -8458 317574
rect -8374 317338 -8138 317574
rect -8694 281658 -8458 281894
rect -8374 281658 -8138 281894
rect -8694 281338 -8458 281574
rect -8374 281338 -8138 281574
rect -8694 245658 -8458 245894
rect -8374 245658 -8138 245894
rect -8694 245338 -8458 245574
rect -8374 245338 -8138 245574
rect -8694 209658 -8458 209894
rect -8374 209658 -8138 209894
rect -8694 209338 -8458 209574
rect -8374 209338 -8138 209574
rect -8694 173658 -8458 173894
rect -8374 173658 -8138 173894
rect -8694 173338 -8458 173574
rect -8374 173338 -8138 173574
rect -8694 137658 -8458 137894
rect -8374 137658 -8138 137894
rect -8694 137338 -8458 137574
rect -8374 137338 -8138 137574
rect -8694 101658 -8458 101894
rect -8374 101658 -8138 101894
rect -8694 101338 -8458 101574
rect -8374 101338 -8138 101574
rect -8694 65658 -8458 65894
rect -8374 65658 -8138 65894
rect -8694 65338 -8458 65574
rect -8374 65338 -8138 65574
rect -8694 29658 -8458 29894
rect -8374 29658 -8138 29894
rect -8694 29338 -8458 29574
rect -8374 29338 -8138 29574
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673938 -7498 674174
rect -7414 673938 -7178 674174
rect -7734 673618 -7498 673854
rect -7414 673618 -7178 673854
rect -7734 637938 -7498 638174
rect -7414 637938 -7178 638174
rect -7734 637618 -7498 637854
rect -7414 637618 -7178 637854
rect -7734 601938 -7498 602174
rect -7414 601938 -7178 602174
rect -7734 601618 -7498 601854
rect -7414 601618 -7178 601854
rect -7734 565938 -7498 566174
rect -7414 565938 -7178 566174
rect -7734 565618 -7498 565854
rect -7414 565618 -7178 565854
rect -7734 529938 -7498 530174
rect -7414 529938 -7178 530174
rect -7734 529618 -7498 529854
rect -7414 529618 -7178 529854
rect -7734 493938 -7498 494174
rect -7414 493938 -7178 494174
rect -7734 493618 -7498 493854
rect -7414 493618 -7178 493854
rect -7734 457938 -7498 458174
rect -7414 457938 -7178 458174
rect -7734 457618 -7498 457854
rect -7414 457618 -7178 457854
rect -7734 421938 -7498 422174
rect -7414 421938 -7178 422174
rect -7734 421618 -7498 421854
rect -7414 421618 -7178 421854
rect -7734 385938 -7498 386174
rect -7414 385938 -7178 386174
rect -7734 385618 -7498 385854
rect -7414 385618 -7178 385854
rect -7734 349938 -7498 350174
rect -7414 349938 -7178 350174
rect -7734 349618 -7498 349854
rect -7414 349618 -7178 349854
rect -7734 313938 -7498 314174
rect -7414 313938 -7178 314174
rect -7734 313618 -7498 313854
rect -7414 313618 -7178 313854
rect -7734 277938 -7498 278174
rect -7414 277938 -7178 278174
rect -7734 277618 -7498 277854
rect -7414 277618 -7178 277854
rect -7734 241938 -7498 242174
rect -7414 241938 -7178 242174
rect -7734 241618 -7498 241854
rect -7414 241618 -7178 241854
rect -7734 205938 -7498 206174
rect -7414 205938 -7178 206174
rect -7734 205618 -7498 205854
rect -7414 205618 -7178 205854
rect -7734 169938 -7498 170174
rect -7414 169938 -7178 170174
rect -7734 169618 -7498 169854
rect -7414 169618 -7178 169854
rect -7734 133938 -7498 134174
rect -7414 133938 -7178 134174
rect -7734 133618 -7498 133854
rect -7414 133618 -7178 133854
rect -7734 97938 -7498 98174
rect -7414 97938 -7178 98174
rect -7734 97618 -7498 97854
rect -7414 97618 -7178 97854
rect -7734 61938 -7498 62174
rect -7414 61938 -7178 62174
rect -7734 61618 -7498 61854
rect -7414 61618 -7178 61854
rect -7734 25938 -7498 26174
rect -7414 25938 -7178 26174
rect -7734 25618 -7498 25854
rect -7414 25618 -7178 25854
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 670218 -6538 670454
rect -6454 670218 -6218 670454
rect -6774 669898 -6538 670134
rect -6454 669898 -6218 670134
rect -6774 634218 -6538 634454
rect -6454 634218 -6218 634454
rect -6774 633898 -6538 634134
rect -6454 633898 -6218 634134
rect -6774 598218 -6538 598454
rect -6454 598218 -6218 598454
rect -6774 597898 -6538 598134
rect -6454 597898 -6218 598134
rect -6774 562218 -6538 562454
rect -6454 562218 -6218 562454
rect -6774 561898 -6538 562134
rect -6454 561898 -6218 562134
rect -6774 526218 -6538 526454
rect -6454 526218 -6218 526454
rect -6774 525898 -6538 526134
rect -6454 525898 -6218 526134
rect -6774 490218 -6538 490454
rect -6454 490218 -6218 490454
rect -6774 489898 -6538 490134
rect -6454 489898 -6218 490134
rect -6774 454218 -6538 454454
rect -6454 454218 -6218 454454
rect -6774 453898 -6538 454134
rect -6454 453898 -6218 454134
rect -6774 418218 -6538 418454
rect -6454 418218 -6218 418454
rect -6774 417898 -6538 418134
rect -6454 417898 -6218 418134
rect -6774 382218 -6538 382454
rect -6454 382218 -6218 382454
rect -6774 381898 -6538 382134
rect -6454 381898 -6218 382134
rect -6774 346218 -6538 346454
rect -6454 346218 -6218 346454
rect -6774 345898 -6538 346134
rect -6454 345898 -6218 346134
rect -6774 310218 -6538 310454
rect -6454 310218 -6218 310454
rect -6774 309898 -6538 310134
rect -6454 309898 -6218 310134
rect -6774 274218 -6538 274454
rect -6454 274218 -6218 274454
rect -6774 273898 -6538 274134
rect -6454 273898 -6218 274134
rect -6774 238218 -6538 238454
rect -6454 238218 -6218 238454
rect -6774 237898 -6538 238134
rect -6454 237898 -6218 238134
rect -6774 202218 -6538 202454
rect -6454 202218 -6218 202454
rect -6774 201898 -6538 202134
rect -6454 201898 -6218 202134
rect -6774 166218 -6538 166454
rect -6454 166218 -6218 166454
rect -6774 165898 -6538 166134
rect -6454 165898 -6218 166134
rect -6774 130218 -6538 130454
rect -6454 130218 -6218 130454
rect -6774 129898 -6538 130134
rect -6454 129898 -6218 130134
rect -6774 94218 -6538 94454
rect -6454 94218 -6218 94454
rect -6774 93898 -6538 94134
rect -6454 93898 -6218 94134
rect -6774 58218 -6538 58454
rect -6454 58218 -6218 58454
rect -6774 57898 -6538 58134
rect -6454 57898 -6218 58134
rect -6774 22218 -6538 22454
rect -6454 22218 -6218 22454
rect -6774 21898 -6538 22134
rect -6454 21898 -6218 22134
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666498 -5578 666734
rect -5494 666498 -5258 666734
rect -5814 666178 -5578 666414
rect -5494 666178 -5258 666414
rect -5814 630498 -5578 630734
rect -5494 630498 -5258 630734
rect -5814 630178 -5578 630414
rect -5494 630178 -5258 630414
rect -5814 594498 -5578 594734
rect -5494 594498 -5258 594734
rect -5814 594178 -5578 594414
rect -5494 594178 -5258 594414
rect -5814 558498 -5578 558734
rect -5494 558498 -5258 558734
rect -5814 558178 -5578 558414
rect -5494 558178 -5258 558414
rect -5814 522498 -5578 522734
rect -5494 522498 -5258 522734
rect -5814 522178 -5578 522414
rect -5494 522178 -5258 522414
rect -5814 486498 -5578 486734
rect -5494 486498 -5258 486734
rect -5814 486178 -5578 486414
rect -5494 486178 -5258 486414
rect -5814 450498 -5578 450734
rect -5494 450498 -5258 450734
rect -5814 450178 -5578 450414
rect -5494 450178 -5258 450414
rect -5814 414498 -5578 414734
rect -5494 414498 -5258 414734
rect -5814 414178 -5578 414414
rect -5494 414178 -5258 414414
rect -5814 378498 -5578 378734
rect -5494 378498 -5258 378734
rect -5814 378178 -5578 378414
rect -5494 378178 -5258 378414
rect -5814 342498 -5578 342734
rect -5494 342498 -5258 342734
rect -5814 342178 -5578 342414
rect -5494 342178 -5258 342414
rect -5814 306498 -5578 306734
rect -5494 306498 -5258 306734
rect -5814 306178 -5578 306414
rect -5494 306178 -5258 306414
rect -5814 270498 -5578 270734
rect -5494 270498 -5258 270734
rect -5814 270178 -5578 270414
rect -5494 270178 -5258 270414
rect -5814 234498 -5578 234734
rect -5494 234498 -5258 234734
rect -5814 234178 -5578 234414
rect -5494 234178 -5258 234414
rect -5814 198498 -5578 198734
rect -5494 198498 -5258 198734
rect -5814 198178 -5578 198414
rect -5494 198178 -5258 198414
rect -5814 162498 -5578 162734
rect -5494 162498 -5258 162734
rect -5814 162178 -5578 162414
rect -5494 162178 -5258 162414
rect -5814 126498 -5578 126734
rect -5494 126498 -5258 126734
rect -5814 126178 -5578 126414
rect -5494 126178 -5258 126414
rect -5814 90498 -5578 90734
rect -5494 90498 -5258 90734
rect -5814 90178 -5578 90414
rect -5494 90178 -5258 90414
rect -5814 54498 -5578 54734
rect -5494 54498 -5258 54734
rect -5814 54178 -5578 54414
rect -5494 54178 -5258 54414
rect -5814 18498 -5578 18734
rect -5494 18498 -5258 18734
rect -5814 18178 -5578 18414
rect -5494 18178 -5258 18414
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698778 -4618 699014
rect -4534 698778 -4298 699014
rect -4854 698458 -4618 698694
rect -4534 698458 -4298 698694
rect -4854 662778 -4618 663014
rect -4534 662778 -4298 663014
rect -4854 662458 -4618 662694
rect -4534 662458 -4298 662694
rect -4854 626778 -4618 627014
rect -4534 626778 -4298 627014
rect -4854 626458 -4618 626694
rect -4534 626458 -4298 626694
rect -4854 590778 -4618 591014
rect -4534 590778 -4298 591014
rect -4854 590458 -4618 590694
rect -4534 590458 -4298 590694
rect -4854 554778 -4618 555014
rect -4534 554778 -4298 555014
rect -4854 554458 -4618 554694
rect -4534 554458 -4298 554694
rect -4854 518778 -4618 519014
rect -4534 518778 -4298 519014
rect -4854 518458 -4618 518694
rect -4534 518458 -4298 518694
rect -4854 482778 -4618 483014
rect -4534 482778 -4298 483014
rect -4854 482458 -4618 482694
rect -4534 482458 -4298 482694
rect -4854 446778 -4618 447014
rect -4534 446778 -4298 447014
rect -4854 446458 -4618 446694
rect -4534 446458 -4298 446694
rect -4854 410778 -4618 411014
rect -4534 410778 -4298 411014
rect -4854 410458 -4618 410694
rect -4534 410458 -4298 410694
rect -4854 374778 -4618 375014
rect -4534 374778 -4298 375014
rect -4854 374458 -4618 374694
rect -4534 374458 -4298 374694
rect -4854 338778 -4618 339014
rect -4534 338778 -4298 339014
rect -4854 338458 -4618 338694
rect -4534 338458 -4298 338694
rect -4854 302778 -4618 303014
rect -4534 302778 -4298 303014
rect -4854 302458 -4618 302694
rect -4534 302458 -4298 302694
rect -4854 266778 -4618 267014
rect -4534 266778 -4298 267014
rect -4854 266458 -4618 266694
rect -4534 266458 -4298 266694
rect -4854 230778 -4618 231014
rect -4534 230778 -4298 231014
rect -4854 230458 -4618 230694
rect -4534 230458 -4298 230694
rect -4854 194778 -4618 195014
rect -4534 194778 -4298 195014
rect -4854 194458 -4618 194694
rect -4534 194458 -4298 194694
rect -4854 158778 -4618 159014
rect -4534 158778 -4298 159014
rect -4854 158458 -4618 158694
rect -4534 158458 -4298 158694
rect -4854 122778 -4618 123014
rect -4534 122778 -4298 123014
rect -4854 122458 -4618 122694
rect -4534 122458 -4298 122694
rect -4854 86778 -4618 87014
rect -4534 86778 -4298 87014
rect -4854 86458 -4618 86694
rect -4534 86458 -4298 86694
rect -4854 50778 -4618 51014
rect -4534 50778 -4298 51014
rect -4854 50458 -4618 50694
rect -4534 50458 -4298 50694
rect -4854 14778 -4618 15014
rect -4534 14778 -4298 15014
rect -4854 14458 -4618 14694
rect -4534 14458 -4298 14694
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 695058 -3658 695294
rect -3574 695058 -3338 695294
rect -3894 694738 -3658 694974
rect -3574 694738 -3338 694974
rect -3894 659058 -3658 659294
rect -3574 659058 -3338 659294
rect -3894 658738 -3658 658974
rect -3574 658738 -3338 658974
rect -3894 623058 -3658 623294
rect -3574 623058 -3338 623294
rect -3894 622738 -3658 622974
rect -3574 622738 -3338 622974
rect -3894 587058 -3658 587294
rect -3574 587058 -3338 587294
rect -3894 586738 -3658 586974
rect -3574 586738 -3338 586974
rect -3894 551058 -3658 551294
rect -3574 551058 -3338 551294
rect -3894 550738 -3658 550974
rect -3574 550738 -3338 550974
rect -3894 515058 -3658 515294
rect -3574 515058 -3338 515294
rect -3894 514738 -3658 514974
rect -3574 514738 -3338 514974
rect -3894 479058 -3658 479294
rect -3574 479058 -3338 479294
rect -3894 478738 -3658 478974
rect -3574 478738 -3338 478974
rect -3894 443058 -3658 443294
rect -3574 443058 -3338 443294
rect -3894 442738 -3658 442974
rect -3574 442738 -3338 442974
rect -3894 407058 -3658 407294
rect -3574 407058 -3338 407294
rect -3894 406738 -3658 406974
rect -3574 406738 -3338 406974
rect -3894 371058 -3658 371294
rect -3574 371058 -3338 371294
rect -3894 370738 -3658 370974
rect -3574 370738 -3338 370974
rect -3894 335058 -3658 335294
rect -3574 335058 -3338 335294
rect -3894 334738 -3658 334974
rect -3574 334738 -3338 334974
rect -3894 299058 -3658 299294
rect -3574 299058 -3338 299294
rect -3894 298738 -3658 298974
rect -3574 298738 -3338 298974
rect -3894 263058 -3658 263294
rect -3574 263058 -3338 263294
rect -3894 262738 -3658 262974
rect -3574 262738 -3338 262974
rect -3894 227058 -3658 227294
rect -3574 227058 -3338 227294
rect -3894 226738 -3658 226974
rect -3574 226738 -3338 226974
rect -3894 191058 -3658 191294
rect -3574 191058 -3338 191294
rect -3894 190738 -3658 190974
rect -3574 190738 -3338 190974
rect -3894 155058 -3658 155294
rect -3574 155058 -3338 155294
rect -3894 154738 -3658 154974
rect -3574 154738 -3338 154974
rect -3894 119058 -3658 119294
rect -3574 119058 -3338 119294
rect -3894 118738 -3658 118974
rect -3574 118738 -3338 118974
rect -3894 83058 -3658 83294
rect -3574 83058 -3338 83294
rect -3894 82738 -3658 82974
rect -3574 82738 -3338 82974
rect -3894 47058 -3658 47294
rect -3574 47058 -3338 47294
rect -3894 46738 -3658 46974
rect -3574 46738 -3338 46974
rect -3894 11058 -3658 11294
rect -3574 11058 -3338 11294
rect -3894 10738 -3658 10974
rect -3574 10738 -3338 10974
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691338 -2698 691574
rect -2614 691338 -2378 691574
rect -2934 691018 -2698 691254
rect -2614 691018 -2378 691254
rect -2934 655338 -2698 655574
rect -2614 655338 -2378 655574
rect -2934 655018 -2698 655254
rect -2614 655018 -2378 655254
rect -2934 619338 -2698 619574
rect -2614 619338 -2378 619574
rect -2934 619018 -2698 619254
rect -2614 619018 -2378 619254
rect -2934 583338 -2698 583574
rect -2614 583338 -2378 583574
rect -2934 583018 -2698 583254
rect -2614 583018 -2378 583254
rect -2934 547338 -2698 547574
rect -2614 547338 -2378 547574
rect -2934 547018 -2698 547254
rect -2614 547018 -2378 547254
rect -2934 511338 -2698 511574
rect -2614 511338 -2378 511574
rect -2934 511018 -2698 511254
rect -2614 511018 -2378 511254
rect -2934 475338 -2698 475574
rect -2614 475338 -2378 475574
rect -2934 475018 -2698 475254
rect -2614 475018 -2378 475254
rect -2934 439338 -2698 439574
rect -2614 439338 -2378 439574
rect -2934 439018 -2698 439254
rect -2614 439018 -2378 439254
rect -2934 403338 -2698 403574
rect -2614 403338 -2378 403574
rect -2934 403018 -2698 403254
rect -2614 403018 -2378 403254
rect -2934 367338 -2698 367574
rect -2614 367338 -2378 367574
rect -2934 367018 -2698 367254
rect -2614 367018 -2378 367254
rect -2934 331338 -2698 331574
rect -2614 331338 -2378 331574
rect -2934 331018 -2698 331254
rect -2614 331018 -2378 331254
rect -2934 295338 -2698 295574
rect -2614 295338 -2378 295574
rect -2934 295018 -2698 295254
rect -2614 295018 -2378 295254
rect -2934 259338 -2698 259574
rect -2614 259338 -2378 259574
rect -2934 259018 -2698 259254
rect -2614 259018 -2378 259254
rect -2934 223338 -2698 223574
rect -2614 223338 -2378 223574
rect -2934 223018 -2698 223254
rect -2614 223018 -2378 223254
rect -2934 187338 -2698 187574
rect -2614 187338 -2378 187574
rect -2934 187018 -2698 187254
rect -2614 187018 -2378 187254
rect -2934 151338 -2698 151574
rect -2614 151338 -2378 151574
rect -2934 151018 -2698 151254
rect -2614 151018 -2378 151254
rect -2934 115338 -2698 115574
rect -2614 115338 -2378 115574
rect -2934 115018 -2698 115254
rect -2614 115018 -2378 115254
rect -2934 79338 -2698 79574
rect -2614 79338 -2378 79574
rect -2934 79018 -2698 79254
rect -2614 79018 -2378 79254
rect -2934 43338 -2698 43574
rect -2614 43338 -2378 43574
rect -2934 43018 -2698 43254
rect -2614 43018 -2378 43254
rect -2934 7338 -2698 7574
rect -2614 7338 -2378 7574
rect -2934 7018 -2698 7254
rect -2614 7018 -2378 7254
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687618 -1738 687854
rect -1654 687618 -1418 687854
rect -1974 687298 -1738 687534
rect -1654 687298 -1418 687534
rect -1974 651618 -1738 651854
rect -1654 651618 -1418 651854
rect -1974 651298 -1738 651534
rect -1654 651298 -1418 651534
rect -1974 615618 -1738 615854
rect -1654 615618 -1418 615854
rect -1974 615298 -1738 615534
rect -1654 615298 -1418 615534
rect -1974 579618 -1738 579854
rect -1654 579618 -1418 579854
rect -1974 579298 -1738 579534
rect -1654 579298 -1418 579534
rect -1974 543618 -1738 543854
rect -1654 543618 -1418 543854
rect -1974 543298 -1738 543534
rect -1654 543298 -1418 543534
rect -1974 507618 -1738 507854
rect -1654 507618 -1418 507854
rect -1974 507298 -1738 507534
rect -1654 507298 -1418 507534
rect -1974 471618 -1738 471854
rect -1654 471618 -1418 471854
rect -1974 471298 -1738 471534
rect -1654 471298 -1418 471534
rect -1974 435618 -1738 435854
rect -1654 435618 -1418 435854
rect -1974 435298 -1738 435534
rect -1654 435298 -1418 435534
rect -1974 399618 -1738 399854
rect -1654 399618 -1418 399854
rect -1974 399298 -1738 399534
rect -1654 399298 -1418 399534
rect -1974 363618 -1738 363854
rect -1654 363618 -1418 363854
rect -1974 363298 -1738 363534
rect -1654 363298 -1418 363534
rect -1974 327618 -1738 327854
rect -1654 327618 -1418 327854
rect -1974 327298 -1738 327534
rect -1654 327298 -1418 327534
rect -1974 291618 -1738 291854
rect -1654 291618 -1418 291854
rect -1974 291298 -1738 291534
rect -1654 291298 -1418 291534
rect -1974 255618 -1738 255854
rect -1654 255618 -1418 255854
rect -1974 255298 -1738 255534
rect -1654 255298 -1418 255534
rect -1974 219618 -1738 219854
rect -1654 219618 -1418 219854
rect -1974 219298 -1738 219534
rect -1654 219298 -1418 219534
rect -1974 183618 -1738 183854
rect -1654 183618 -1418 183854
rect -1974 183298 -1738 183534
rect -1654 183298 -1418 183534
rect -1974 147618 -1738 147854
rect -1654 147618 -1418 147854
rect -1974 147298 -1738 147534
rect -1654 147298 -1418 147534
rect -1974 111618 -1738 111854
rect -1654 111618 -1418 111854
rect -1974 111298 -1738 111534
rect -1654 111298 -1418 111534
rect -1974 75618 -1738 75854
rect -1654 75618 -1418 75854
rect -1974 75298 -1738 75534
rect -1654 75298 -1418 75534
rect -1974 39618 -1738 39854
rect -1654 39618 -1418 39854
rect -1974 39298 -1738 39534
rect -1654 39298 -1418 39534
rect -1974 3618 -1738 3854
rect -1654 3618 -1418 3854
rect -1974 3298 -1738 3534
rect -1654 3298 -1418 3534
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 2226 704602 2462 704838
rect 2546 704602 2782 704838
rect 2226 704282 2462 704518
rect 2546 704282 2782 704518
rect 2226 687618 2462 687854
rect 2546 687618 2782 687854
rect 2226 687298 2462 687534
rect 2546 687298 2782 687534
rect 2226 651618 2462 651854
rect 2546 651618 2782 651854
rect 2226 651298 2462 651534
rect 2546 651298 2782 651534
rect 2226 615618 2462 615854
rect 2546 615618 2782 615854
rect 2226 615298 2462 615534
rect 2546 615298 2782 615534
rect 2226 579618 2462 579854
rect 2546 579618 2782 579854
rect 2226 579298 2462 579534
rect 2546 579298 2782 579534
rect 2226 543618 2462 543854
rect 2546 543618 2782 543854
rect 2226 543298 2462 543534
rect 2546 543298 2782 543534
rect 2226 507618 2462 507854
rect 2546 507618 2782 507854
rect 2226 507298 2462 507534
rect 2546 507298 2782 507534
rect 2226 471618 2462 471854
rect 2546 471618 2782 471854
rect 2226 471298 2462 471534
rect 2546 471298 2782 471534
rect 2226 435618 2462 435854
rect 2546 435618 2782 435854
rect 2226 435298 2462 435534
rect 2546 435298 2782 435534
rect 2226 399618 2462 399854
rect 2546 399618 2782 399854
rect 2226 399298 2462 399534
rect 2546 399298 2782 399534
rect 2226 363618 2462 363854
rect 2546 363618 2782 363854
rect 2226 363298 2462 363534
rect 2546 363298 2782 363534
rect 2226 327618 2462 327854
rect 2546 327618 2782 327854
rect 2226 327298 2462 327534
rect 2546 327298 2782 327534
rect 2226 291618 2462 291854
rect 2546 291618 2782 291854
rect 2226 291298 2462 291534
rect 2546 291298 2782 291534
rect 2226 255618 2462 255854
rect 2546 255618 2782 255854
rect 2226 255298 2462 255534
rect 2546 255298 2782 255534
rect 2226 219618 2462 219854
rect 2546 219618 2782 219854
rect 2226 219298 2462 219534
rect 2546 219298 2782 219534
rect 2226 183618 2462 183854
rect 2546 183618 2782 183854
rect 2226 183298 2462 183534
rect 2546 183298 2782 183534
rect 2226 147618 2462 147854
rect 2546 147618 2782 147854
rect 2226 147298 2462 147534
rect 2546 147298 2782 147534
rect 2226 111618 2462 111854
rect 2546 111618 2782 111854
rect 2226 111298 2462 111534
rect 2546 111298 2782 111534
rect 2226 75618 2462 75854
rect 2546 75618 2782 75854
rect 2226 75298 2462 75534
rect 2546 75298 2782 75534
rect 2226 39618 2462 39854
rect 2546 39618 2782 39854
rect 2226 39298 2462 39534
rect 2546 39298 2782 39534
rect 2226 3618 2462 3854
rect 2546 3618 2782 3854
rect 2226 3298 2462 3534
rect 2546 3298 2782 3534
rect 2226 -582 2462 -346
rect 2546 -582 2782 -346
rect 2226 -902 2462 -666
rect 2546 -902 2782 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5946 705562 6182 705798
rect 6266 705562 6502 705798
rect 5946 705242 6182 705478
rect 6266 705242 6502 705478
rect 5946 691338 6182 691574
rect 6266 691338 6502 691574
rect 5946 691018 6182 691254
rect 6266 691018 6502 691254
rect 5946 655338 6182 655574
rect 6266 655338 6502 655574
rect 5946 655018 6182 655254
rect 6266 655018 6502 655254
rect 5946 619338 6182 619574
rect 6266 619338 6502 619574
rect 5946 619018 6182 619254
rect 6266 619018 6502 619254
rect 5946 583338 6182 583574
rect 6266 583338 6502 583574
rect 5946 583018 6182 583254
rect 6266 583018 6502 583254
rect 5946 547338 6182 547574
rect 6266 547338 6502 547574
rect 5946 547018 6182 547254
rect 6266 547018 6502 547254
rect 5946 511338 6182 511574
rect 6266 511338 6502 511574
rect 5946 511018 6182 511254
rect 6266 511018 6502 511254
rect 5946 475338 6182 475574
rect 6266 475338 6502 475574
rect 5946 475018 6182 475254
rect 6266 475018 6502 475254
rect 5946 439338 6182 439574
rect 6266 439338 6502 439574
rect 5946 439018 6182 439254
rect 6266 439018 6502 439254
rect 5946 403338 6182 403574
rect 6266 403338 6502 403574
rect 5946 403018 6182 403254
rect 6266 403018 6502 403254
rect 5946 367338 6182 367574
rect 6266 367338 6502 367574
rect 5946 367018 6182 367254
rect 6266 367018 6502 367254
rect 5946 331338 6182 331574
rect 6266 331338 6502 331574
rect 5946 331018 6182 331254
rect 6266 331018 6502 331254
rect 5946 295338 6182 295574
rect 6266 295338 6502 295574
rect 5946 295018 6182 295254
rect 6266 295018 6502 295254
rect 5946 259338 6182 259574
rect 6266 259338 6502 259574
rect 5946 259018 6182 259254
rect 6266 259018 6502 259254
rect 5946 223338 6182 223574
rect 6266 223338 6502 223574
rect 5946 223018 6182 223254
rect 6266 223018 6502 223254
rect 5946 187338 6182 187574
rect 6266 187338 6502 187574
rect 5946 187018 6182 187254
rect 6266 187018 6502 187254
rect 5946 151338 6182 151574
rect 6266 151338 6502 151574
rect 5946 151018 6182 151254
rect 6266 151018 6502 151254
rect 5946 115338 6182 115574
rect 6266 115338 6502 115574
rect 5946 115018 6182 115254
rect 6266 115018 6502 115254
rect 5946 79338 6182 79574
rect 6266 79338 6502 79574
rect 5946 79018 6182 79254
rect 6266 79018 6502 79254
rect 5946 43338 6182 43574
rect 6266 43338 6502 43574
rect 5946 43018 6182 43254
rect 6266 43018 6502 43254
rect 5946 7338 6182 7574
rect 6266 7338 6502 7574
rect 5946 7018 6182 7254
rect 6266 7018 6502 7254
rect 5946 -1542 6182 -1306
rect 6266 -1542 6502 -1306
rect 5946 -1862 6182 -1626
rect 6266 -1862 6502 -1626
rect 9666 706522 9902 706758
rect 9986 706522 10222 706758
rect 9666 706202 9902 706438
rect 9986 706202 10222 706438
rect 9666 695058 9902 695294
rect 9986 695058 10222 695294
rect 9666 694738 9902 694974
rect 9986 694738 10222 694974
rect 9666 659058 9902 659294
rect 9986 659058 10222 659294
rect 9666 658738 9902 658974
rect 9986 658738 10222 658974
rect 9666 623058 9902 623294
rect 9986 623058 10222 623294
rect 9666 622738 9902 622974
rect 9986 622738 10222 622974
rect 9666 587058 9902 587294
rect 9986 587058 10222 587294
rect 9666 586738 9902 586974
rect 9986 586738 10222 586974
rect 9666 551058 9902 551294
rect 9986 551058 10222 551294
rect 9666 550738 9902 550974
rect 9986 550738 10222 550974
rect 9666 515058 9902 515294
rect 9986 515058 10222 515294
rect 9666 514738 9902 514974
rect 9986 514738 10222 514974
rect 9666 479058 9902 479294
rect 9986 479058 10222 479294
rect 9666 478738 9902 478974
rect 9986 478738 10222 478974
rect 9666 443058 9902 443294
rect 9986 443058 10222 443294
rect 9666 442738 9902 442974
rect 9986 442738 10222 442974
rect 9666 407058 9902 407294
rect 9986 407058 10222 407294
rect 9666 406738 9902 406974
rect 9986 406738 10222 406974
rect 9666 371058 9902 371294
rect 9986 371058 10222 371294
rect 9666 370738 9902 370974
rect 9986 370738 10222 370974
rect 9666 335058 9902 335294
rect 9986 335058 10222 335294
rect 9666 334738 9902 334974
rect 9986 334738 10222 334974
rect 9666 299058 9902 299294
rect 9986 299058 10222 299294
rect 9666 298738 9902 298974
rect 9986 298738 10222 298974
rect 9666 263058 9902 263294
rect 9986 263058 10222 263294
rect 9666 262738 9902 262974
rect 9986 262738 10222 262974
rect 9666 227058 9902 227294
rect 9986 227058 10222 227294
rect 9666 226738 9902 226974
rect 9986 226738 10222 226974
rect 9666 191058 9902 191294
rect 9986 191058 10222 191294
rect 9666 190738 9902 190974
rect 9986 190738 10222 190974
rect 9666 155058 9902 155294
rect 9986 155058 10222 155294
rect 9666 154738 9902 154974
rect 9986 154738 10222 154974
rect 9666 119058 9902 119294
rect 9986 119058 10222 119294
rect 9666 118738 9902 118974
rect 9986 118738 10222 118974
rect 9666 83058 9902 83294
rect 9986 83058 10222 83294
rect 9666 82738 9902 82974
rect 9986 82738 10222 82974
rect 9666 47058 9902 47294
rect 9986 47058 10222 47294
rect 9666 46738 9902 46974
rect 9986 46738 10222 46974
rect 9666 11058 9902 11294
rect 9986 11058 10222 11294
rect 9666 10738 9902 10974
rect 9986 10738 10222 10974
rect 13386 707482 13622 707718
rect 13706 707482 13942 707718
rect 13386 707162 13622 707398
rect 13706 707162 13942 707398
rect 13386 698778 13622 699014
rect 13706 698778 13942 699014
rect 13386 698458 13622 698694
rect 13706 698458 13942 698694
rect 13386 662778 13622 663014
rect 13706 662778 13942 663014
rect 13386 662458 13622 662694
rect 13706 662458 13942 662694
rect 13386 626778 13622 627014
rect 13706 626778 13942 627014
rect 13386 626458 13622 626694
rect 13706 626458 13942 626694
rect 13386 590778 13622 591014
rect 13706 590778 13942 591014
rect 13386 590458 13622 590694
rect 13706 590458 13942 590694
rect 13386 554778 13622 555014
rect 13706 554778 13942 555014
rect 13386 554458 13622 554694
rect 13706 554458 13942 554694
rect 13386 518778 13622 519014
rect 13706 518778 13942 519014
rect 13386 518458 13622 518694
rect 13706 518458 13942 518694
rect 13386 482778 13622 483014
rect 13706 482778 13942 483014
rect 13386 482458 13622 482694
rect 13706 482458 13942 482694
rect 13386 446778 13622 447014
rect 13706 446778 13942 447014
rect 13386 446458 13622 446694
rect 13706 446458 13942 446694
rect 13386 410778 13622 411014
rect 13706 410778 13942 411014
rect 13386 410458 13622 410694
rect 13706 410458 13942 410694
rect 13386 374778 13622 375014
rect 13706 374778 13942 375014
rect 13386 374458 13622 374694
rect 13706 374458 13942 374694
rect 13386 338778 13622 339014
rect 13706 338778 13942 339014
rect 13386 338458 13622 338694
rect 13706 338458 13942 338694
rect 13386 302778 13622 303014
rect 13706 302778 13942 303014
rect 13386 302458 13622 302694
rect 13706 302458 13942 302694
rect 13386 266778 13622 267014
rect 13706 266778 13942 267014
rect 13386 266458 13622 266694
rect 13706 266458 13942 266694
rect 13386 230778 13622 231014
rect 13706 230778 13942 231014
rect 13386 230458 13622 230694
rect 13706 230458 13942 230694
rect 13386 194778 13622 195014
rect 13706 194778 13942 195014
rect 13386 194458 13622 194694
rect 13706 194458 13942 194694
rect 13386 158778 13622 159014
rect 13706 158778 13942 159014
rect 13386 158458 13622 158694
rect 13706 158458 13942 158694
rect 13386 122778 13622 123014
rect 13706 122778 13942 123014
rect 13386 122458 13622 122694
rect 13706 122458 13942 122694
rect 13386 86778 13622 87014
rect 13706 86778 13942 87014
rect 13386 86458 13622 86694
rect 13706 86458 13942 86694
rect 13386 50778 13622 51014
rect 13706 50778 13942 51014
rect 13386 50458 13622 50694
rect 13706 50458 13942 50694
rect 13386 14778 13622 15014
rect 13706 14778 13942 15014
rect 13386 14458 13622 14694
rect 13706 14458 13942 14694
rect 12302 4302 12538 4538
rect 9666 -2502 9902 -2266
rect 9986 -2502 10222 -2266
rect 9666 -2822 9902 -2586
rect 9986 -2822 10222 -2586
rect 13386 -3462 13622 -3226
rect 13706 -3462 13942 -3226
rect 13386 -3782 13622 -3546
rect 13706 -3782 13942 -3546
rect 17106 708442 17342 708678
rect 17426 708442 17662 708678
rect 17106 708122 17342 708358
rect 17426 708122 17662 708358
rect 17106 666498 17342 666734
rect 17426 666498 17662 666734
rect 17106 666178 17342 666414
rect 17426 666178 17662 666414
rect 17106 630498 17342 630734
rect 17426 630498 17662 630734
rect 17106 630178 17342 630414
rect 17426 630178 17662 630414
rect 17106 594498 17342 594734
rect 17426 594498 17662 594734
rect 17106 594178 17342 594414
rect 17426 594178 17662 594414
rect 17106 558498 17342 558734
rect 17426 558498 17662 558734
rect 17106 558178 17342 558414
rect 17426 558178 17662 558414
rect 17106 522498 17342 522734
rect 17426 522498 17662 522734
rect 17106 522178 17342 522414
rect 17426 522178 17662 522414
rect 17106 486498 17342 486734
rect 17426 486498 17662 486734
rect 17106 486178 17342 486414
rect 17426 486178 17662 486414
rect 17106 450498 17342 450734
rect 17426 450498 17662 450734
rect 17106 450178 17342 450414
rect 17426 450178 17662 450414
rect 17106 414498 17342 414734
rect 17426 414498 17662 414734
rect 17106 414178 17342 414414
rect 17426 414178 17662 414414
rect 17106 378498 17342 378734
rect 17426 378498 17662 378734
rect 17106 378178 17342 378414
rect 17426 378178 17662 378414
rect 17106 342498 17342 342734
rect 17426 342498 17662 342734
rect 17106 342178 17342 342414
rect 17426 342178 17662 342414
rect 17106 306498 17342 306734
rect 17426 306498 17662 306734
rect 17106 306178 17342 306414
rect 17426 306178 17662 306414
rect 17106 270498 17342 270734
rect 17426 270498 17662 270734
rect 17106 270178 17342 270414
rect 17426 270178 17662 270414
rect 17106 234498 17342 234734
rect 17426 234498 17662 234734
rect 17106 234178 17342 234414
rect 17426 234178 17662 234414
rect 17106 198498 17342 198734
rect 17426 198498 17662 198734
rect 17106 198178 17342 198414
rect 17426 198178 17662 198414
rect 17106 162498 17342 162734
rect 17426 162498 17662 162734
rect 17106 162178 17342 162414
rect 17426 162178 17662 162414
rect 17106 126498 17342 126734
rect 17426 126498 17662 126734
rect 17106 126178 17342 126414
rect 17426 126178 17662 126414
rect 17106 90498 17342 90734
rect 17426 90498 17662 90734
rect 17106 90178 17342 90414
rect 17426 90178 17662 90414
rect 17106 54498 17342 54734
rect 17426 54498 17662 54734
rect 17106 54178 17342 54414
rect 17426 54178 17662 54414
rect 17106 18498 17342 18734
rect 17426 18498 17662 18734
rect 17106 18178 17342 18414
rect 17426 18178 17662 18414
rect 17106 -4422 17342 -4186
rect 17426 -4422 17662 -4186
rect 17106 -4742 17342 -4506
rect 17426 -4742 17662 -4506
rect 20826 709402 21062 709638
rect 21146 709402 21382 709638
rect 20826 709082 21062 709318
rect 21146 709082 21382 709318
rect 20826 670218 21062 670454
rect 21146 670218 21382 670454
rect 20826 669898 21062 670134
rect 21146 669898 21382 670134
rect 20826 634218 21062 634454
rect 21146 634218 21382 634454
rect 20826 633898 21062 634134
rect 21146 633898 21382 634134
rect 20826 598218 21062 598454
rect 21146 598218 21382 598454
rect 20826 597898 21062 598134
rect 21146 597898 21382 598134
rect 20826 562218 21062 562454
rect 21146 562218 21382 562454
rect 20826 561898 21062 562134
rect 21146 561898 21382 562134
rect 20826 526218 21062 526454
rect 21146 526218 21382 526454
rect 20826 525898 21062 526134
rect 21146 525898 21382 526134
rect 20826 490218 21062 490454
rect 21146 490218 21382 490454
rect 20826 489898 21062 490134
rect 21146 489898 21382 490134
rect 20826 454218 21062 454454
rect 21146 454218 21382 454454
rect 20826 453898 21062 454134
rect 21146 453898 21382 454134
rect 20826 418218 21062 418454
rect 21146 418218 21382 418454
rect 20826 417898 21062 418134
rect 21146 417898 21382 418134
rect 20826 382218 21062 382454
rect 21146 382218 21382 382454
rect 20826 381898 21062 382134
rect 21146 381898 21382 382134
rect 20826 346218 21062 346454
rect 21146 346218 21382 346454
rect 20826 345898 21062 346134
rect 21146 345898 21382 346134
rect 20826 310218 21062 310454
rect 21146 310218 21382 310454
rect 20826 309898 21062 310134
rect 21146 309898 21382 310134
rect 20826 274218 21062 274454
rect 21146 274218 21382 274454
rect 20826 273898 21062 274134
rect 21146 273898 21382 274134
rect 20826 238218 21062 238454
rect 21146 238218 21382 238454
rect 20826 237898 21062 238134
rect 21146 237898 21382 238134
rect 20826 202218 21062 202454
rect 21146 202218 21382 202454
rect 20826 201898 21062 202134
rect 21146 201898 21382 202134
rect 20826 166218 21062 166454
rect 21146 166218 21382 166454
rect 20826 165898 21062 166134
rect 21146 165898 21382 166134
rect 20826 130218 21062 130454
rect 21146 130218 21382 130454
rect 20826 129898 21062 130134
rect 21146 129898 21382 130134
rect 20826 94218 21062 94454
rect 21146 94218 21382 94454
rect 20826 93898 21062 94134
rect 21146 93898 21382 94134
rect 20826 58218 21062 58454
rect 21146 58218 21382 58454
rect 20826 57898 21062 58134
rect 21146 57898 21382 58134
rect 20826 22218 21062 22454
rect 21146 22218 21382 22454
rect 20826 21898 21062 22134
rect 21146 21898 21382 22134
rect 20826 -5382 21062 -5146
rect 21146 -5382 21382 -5146
rect 20826 -5702 21062 -5466
rect 21146 -5702 21382 -5466
rect 24546 710362 24782 710598
rect 24866 710362 25102 710598
rect 24546 710042 24782 710278
rect 24866 710042 25102 710278
rect 24546 673938 24782 674174
rect 24866 673938 25102 674174
rect 24546 673618 24782 673854
rect 24866 673618 25102 673854
rect 24546 637938 24782 638174
rect 24866 637938 25102 638174
rect 24546 637618 24782 637854
rect 24866 637618 25102 637854
rect 24546 601938 24782 602174
rect 24866 601938 25102 602174
rect 24546 601618 24782 601854
rect 24866 601618 25102 601854
rect 24546 565938 24782 566174
rect 24866 565938 25102 566174
rect 24546 565618 24782 565854
rect 24866 565618 25102 565854
rect 24546 529938 24782 530174
rect 24866 529938 25102 530174
rect 24546 529618 24782 529854
rect 24866 529618 25102 529854
rect 24546 493938 24782 494174
rect 24866 493938 25102 494174
rect 24546 493618 24782 493854
rect 24866 493618 25102 493854
rect 24546 457938 24782 458174
rect 24866 457938 25102 458174
rect 24546 457618 24782 457854
rect 24866 457618 25102 457854
rect 24546 421938 24782 422174
rect 24866 421938 25102 422174
rect 24546 421618 24782 421854
rect 24866 421618 25102 421854
rect 24546 385938 24782 386174
rect 24866 385938 25102 386174
rect 24546 385618 24782 385854
rect 24866 385618 25102 385854
rect 24546 349938 24782 350174
rect 24866 349938 25102 350174
rect 24546 349618 24782 349854
rect 24866 349618 25102 349854
rect 24546 313938 24782 314174
rect 24866 313938 25102 314174
rect 24546 313618 24782 313854
rect 24866 313618 25102 313854
rect 24546 277938 24782 278174
rect 24866 277938 25102 278174
rect 24546 277618 24782 277854
rect 24866 277618 25102 277854
rect 24546 241938 24782 242174
rect 24866 241938 25102 242174
rect 24546 241618 24782 241854
rect 24866 241618 25102 241854
rect 24546 205938 24782 206174
rect 24866 205938 25102 206174
rect 24546 205618 24782 205854
rect 24866 205618 25102 205854
rect 24546 169938 24782 170174
rect 24866 169938 25102 170174
rect 24546 169618 24782 169854
rect 24866 169618 25102 169854
rect 24546 133938 24782 134174
rect 24866 133938 25102 134174
rect 24546 133618 24782 133854
rect 24866 133618 25102 133854
rect 24546 97938 24782 98174
rect 24866 97938 25102 98174
rect 24546 97618 24782 97854
rect 24866 97618 25102 97854
rect 24546 61938 24782 62174
rect 24866 61938 25102 62174
rect 24546 61618 24782 61854
rect 24866 61618 25102 61854
rect 24546 25938 24782 26174
rect 24866 25938 25102 26174
rect 24546 25618 24782 25854
rect 24866 25618 25102 25854
rect 28266 711322 28502 711558
rect 28586 711322 28822 711558
rect 28266 711002 28502 711238
rect 28586 711002 28822 711238
rect 28266 677658 28502 677894
rect 28586 677658 28822 677894
rect 28266 677338 28502 677574
rect 28586 677338 28822 677574
rect 28266 641658 28502 641894
rect 28586 641658 28822 641894
rect 28266 641338 28502 641574
rect 28586 641338 28822 641574
rect 28266 605658 28502 605894
rect 28586 605658 28822 605894
rect 28266 605338 28502 605574
rect 28586 605338 28822 605574
rect 28266 569658 28502 569894
rect 28586 569658 28822 569894
rect 28266 569338 28502 569574
rect 28586 569338 28822 569574
rect 28266 533658 28502 533894
rect 28586 533658 28822 533894
rect 28266 533338 28502 533574
rect 28586 533338 28822 533574
rect 28266 497658 28502 497894
rect 28586 497658 28822 497894
rect 28266 497338 28502 497574
rect 28586 497338 28822 497574
rect 28266 461658 28502 461894
rect 28586 461658 28822 461894
rect 28266 461338 28502 461574
rect 28586 461338 28822 461574
rect 28266 425658 28502 425894
rect 28586 425658 28822 425894
rect 28266 425338 28502 425574
rect 28586 425338 28822 425574
rect 28266 389658 28502 389894
rect 28586 389658 28822 389894
rect 28266 389338 28502 389574
rect 28586 389338 28822 389574
rect 28266 353658 28502 353894
rect 28586 353658 28822 353894
rect 28266 353338 28502 353574
rect 28586 353338 28822 353574
rect 28266 317658 28502 317894
rect 28586 317658 28822 317894
rect 28266 317338 28502 317574
rect 28586 317338 28822 317574
rect 28266 281658 28502 281894
rect 28586 281658 28822 281894
rect 28266 281338 28502 281574
rect 28586 281338 28822 281574
rect 28266 245658 28502 245894
rect 28586 245658 28822 245894
rect 28266 245338 28502 245574
rect 28586 245338 28822 245574
rect 28266 209658 28502 209894
rect 28586 209658 28822 209894
rect 28266 209338 28502 209574
rect 28586 209338 28822 209574
rect 28266 173658 28502 173894
rect 28586 173658 28822 173894
rect 28266 173338 28502 173574
rect 28586 173338 28822 173574
rect 28266 137658 28502 137894
rect 28586 137658 28822 137894
rect 28266 137338 28502 137574
rect 28586 137338 28822 137574
rect 28266 101658 28502 101894
rect 28586 101658 28822 101894
rect 28266 101338 28502 101574
rect 28586 101338 28822 101574
rect 28266 65658 28502 65894
rect 28586 65658 28822 65894
rect 28266 65338 28502 65574
rect 28586 65338 28822 65574
rect 28266 29658 28502 29894
rect 28586 29658 28822 29894
rect 28266 29338 28502 29574
rect 28586 29338 28822 29574
rect 27758 9742 27994 9978
rect 24546 -6342 24782 -6106
rect 24866 -6342 25102 -6106
rect 24546 -6662 24782 -6426
rect 24866 -6662 25102 -6426
rect 28266 -7302 28502 -7066
rect 28586 -7302 28822 -7066
rect 28266 -7622 28502 -7386
rect 28586 -7622 28822 -7386
rect 38226 704602 38462 704838
rect 38546 704602 38782 704838
rect 38226 704282 38462 704518
rect 38546 704282 38782 704518
rect 38226 687618 38462 687854
rect 38546 687618 38782 687854
rect 38226 687298 38462 687534
rect 38546 687298 38782 687534
rect 38226 651618 38462 651854
rect 38546 651618 38782 651854
rect 38226 651298 38462 651534
rect 38546 651298 38782 651534
rect 38226 615618 38462 615854
rect 38546 615618 38782 615854
rect 38226 615298 38462 615534
rect 38546 615298 38782 615534
rect 38226 579618 38462 579854
rect 38546 579618 38782 579854
rect 38226 579298 38462 579534
rect 38546 579298 38782 579534
rect 38226 543618 38462 543854
rect 38546 543618 38782 543854
rect 38226 543298 38462 543534
rect 38546 543298 38782 543534
rect 38226 507618 38462 507854
rect 38546 507618 38782 507854
rect 38226 507298 38462 507534
rect 38546 507298 38782 507534
rect 38226 471618 38462 471854
rect 38546 471618 38782 471854
rect 38226 471298 38462 471534
rect 38546 471298 38782 471534
rect 38226 435618 38462 435854
rect 38546 435618 38782 435854
rect 38226 435298 38462 435534
rect 38546 435298 38782 435534
rect 38226 399618 38462 399854
rect 38546 399618 38782 399854
rect 38226 399298 38462 399534
rect 38546 399298 38782 399534
rect 38226 363618 38462 363854
rect 38546 363618 38782 363854
rect 38226 363298 38462 363534
rect 38546 363298 38782 363534
rect 38226 327618 38462 327854
rect 38546 327618 38782 327854
rect 38226 327298 38462 327534
rect 38546 327298 38782 327534
rect 38226 291618 38462 291854
rect 38546 291618 38782 291854
rect 38226 291298 38462 291534
rect 38546 291298 38782 291534
rect 38226 255618 38462 255854
rect 38546 255618 38782 255854
rect 38226 255298 38462 255534
rect 38546 255298 38782 255534
rect 38226 219618 38462 219854
rect 38546 219618 38782 219854
rect 38226 219298 38462 219534
rect 38546 219298 38782 219534
rect 38226 183618 38462 183854
rect 38546 183618 38782 183854
rect 38226 183298 38462 183534
rect 38546 183298 38782 183534
rect 38226 147618 38462 147854
rect 38546 147618 38782 147854
rect 38226 147298 38462 147534
rect 38546 147298 38782 147534
rect 38226 111618 38462 111854
rect 38546 111618 38782 111854
rect 38226 111298 38462 111534
rect 38546 111298 38782 111534
rect 38226 75618 38462 75854
rect 38546 75618 38782 75854
rect 38226 75298 38462 75534
rect 38546 75298 38782 75534
rect 38226 39618 38462 39854
rect 38546 39618 38782 39854
rect 38226 39298 38462 39534
rect 38546 39298 38782 39534
rect 38226 3618 38462 3854
rect 38546 3618 38782 3854
rect 38226 3298 38462 3534
rect 38546 3298 38782 3534
rect 38226 -582 38462 -346
rect 38546 -582 38782 -346
rect 38226 -902 38462 -666
rect 38546 -902 38782 -666
rect 41946 705562 42182 705798
rect 42266 705562 42502 705798
rect 41946 705242 42182 705478
rect 42266 705242 42502 705478
rect 41946 691338 42182 691574
rect 42266 691338 42502 691574
rect 41946 691018 42182 691254
rect 42266 691018 42502 691254
rect 41946 655338 42182 655574
rect 42266 655338 42502 655574
rect 41946 655018 42182 655254
rect 42266 655018 42502 655254
rect 41946 619338 42182 619574
rect 42266 619338 42502 619574
rect 41946 619018 42182 619254
rect 42266 619018 42502 619254
rect 41946 583338 42182 583574
rect 42266 583338 42502 583574
rect 41946 583018 42182 583254
rect 42266 583018 42502 583254
rect 41946 547338 42182 547574
rect 42266 547338 42502 547574
rect 41946 547018 42182 547254
rect 42266 547018 42502 547254
rect 41946 511338 42182 511574
rect 42266 511338 42502 511574
rect 41946 511018 42182 511254
rect 42266 511018 42502 511254
rect 41946 475338 42182 475574
rect 42266 475338 42502 475574
rect 41946 475018 42182 475254
rect 42266 475018 42502 475254
rect 41946 439338 42182 439574
rect 42266 439338 42502 439574
rect 41946 439018 42182 439254
rect 42266 439018 42502 439254
rect 41946 403338 42182 403574
rect 42266 403338 42502 403574
rect 41946 403018 42182 403254
rect 42266 403018 42502 403254
rect 41946 367338 42182 367574
rect 42266 367338 42502 367574
rect 41946 367018 42182 367254
rect 42266 367018 42502 367254
rect 41946 331338 42182 331574
rect 42266 331338 42502 331574
rect 41946 331018 42182 331254
rect 42266 331018 42502 331254
rect 41946 295338 42182 295574
rect 42266 295338 42502 295574
rect 41946 295018 42182 295254
rect 42266 295018 42502 295254
rect 41946 259338 42182 259574
rect 42266 259338 42502 259574
rect 41946 259018 42182 259254
rect 42266 259018 42502 259254
rect 41946 223338 42182 223574
rect 42266 223338 42502 223574
rect 41946 223018 42182 223254
rect 42266 223018 42502 223254
rect 41946 187338 42182 187574
rect 42266 187338 42502 187574
rect 41946 187018 42182 187254
rect 42266 187018 42502 187254
rect 41946 151338 42182 151574
rect 42266 151338 42502 151574
rect 41946 151018 42182 151254
rect 42266 151018 42502 151254
rect 41946 115338 42182 115574
rect 42266 115338 42502 115574
rect 41946 115018 42182 115254
rect 42266 115018 42502 115254
rect 41946 79338 42182 79574
rect 42266 79338 42502 79574
rect 41946 79018 42182 79254
rect 42266 79018 42502 79254
rect 41946 43338 42182 43574
rect 42266 43338 42502 43574
rect 41946 43018 42182 43254
rect 42266 43018 42502 43254
rect 41946 7338 42182 7574
rect 42266 7338 42502 7574
rect 41946 7018 42182 7254
rect 42266 7018 42502 7254
rect 45666 706522 45902 706758
rect 45986 706522 46222 706758
rect 45666 706202 45902 706438
rect 45986 706202 46222 706438
rect 45666 695058 45902 695294
rect 45986 695058 46222 695294
rect 45666 694738 45902 694974
rect 45986 694738 46222 694974
rect 45666 659058 45902 659294
rect 45986 659058 46222 659294
rect 45666 658738 45902 658974
rect 45986 658738 46222 658974
rect 45666 623058 45902 623294
rect 45986 623058 46222 623294
rect 45666 622738 45902 622974
rect 45986 622738 46222 622974
rect 45666 587058 45902 587294
rect 45986 587058 46222 587294
rect 45666 586738 45902 586974
rect 45986 586738 46222 586974
rect 45666 551058 45902 551294
rect 45986 551058 46222 551294
rect 45666 550738 45902 550974
rect 45986 550738 46222 550974
rect 45666 515058 45902 515294
rect 45986 515058 46222 515294
rect 45666 514738 45902 514974
rect 45986 514738 46222 514974
rect 45666 479058 45902 479294
rect 45986 479058 46222 479294
rect 45666 478738 45902 478974
rect 45986 478738 46222 478974
rect 45666 443058 45902 443294
rect 45986 443058 46222 443294
rect 45666 442738 45902 442974
rect 45986 442738 46222 442974
rect 45666 407058 45902 407294
rect 45986 407058 46222 407294
rect 45666 406738 45902 406974
rect 45986 406738 46222 406974
rect 45666 371058 45902 371294
rect 45986 371058 46222 371294
rect 45666 370738 45902 370974
rect 45986 370738 46222 370974
rect 45666 335058 45902 335294
rect 45986 335058 46222 335294
rect 45666 334738 45902 334974
rect 45986 334738 46222 334974
rect 45666 299058 45902 299294
rect 45986 299058 46222 299294
rect 45666 298738 45902 298974
rect 45986 298738 46222 298974
rect 45666 263058 45902 263294
rect 45986 263058 46222 263294
rect 45666 262738 45902 262974
rect 45986 262738 46222 262974
rect 45666 227058 45902 227294
rect 45986 227058 46222 227294
rect 45666 226738 45902 226974
rect 45986 226738 46222 226974
rect 45666 191058 45902 191294
rect 45986 191058 46222 191294
rect 45666 190738 45902 190974
rect 45986 190738 46222 190974
rect 45666 155058 45902 155294
rect 45986 155058 46222 155294
rect 45666 154738 45902 154974
rect 45986 154738 46222 154974
rect 45666 119058 45902 119294
rect 45986 119058 46222 119294
rect 45666 118738 45902 118974
rect 45986 118738 46222 118974
rect 45666 83058 45902 83294
rect 45986 83058 46222 83294
rect 45666 82738 45902 82974
rect 45986 82738 46222 82974
rect 45666 47058 45902 47294
rect 45986 47058 46222 47294
rect 45666 46738 45902 46974
rect 45986 46738 46222 46974
rect 45666 11058 45902 11294
rect 45986 11058 46222 11294
rect 45666 10738 45902 10974
rect 45986 10738 46222 10974
rect 43950 5662 44186 5898
rect 41946 -1542 42182 -1306
rect 42266 -1542 42502 -1306
rect 41946 -1862 42182 -1626
rect 42266 -1862 42502 -1626
rect 45666 -2502 45902 -2266
rect 45986 -2502 46222 -2266
rect 45666 -2822 45902 -2586
rect 45986 -2822 46222 -2586
rect 49386 707482 49622 707718
rect 49706 707482 49942 707718
rect 49386 707162 49622 707398
rect 49706 707162 49942 707398
rect 49386 698778 49622 699014
rect 49706 698778 49942 699014
rect 49386 698458 49622 698694
rect 49706 698458 49942 698694
rect 49386 662778 49622 663014
rect 49706 662778 49942 663014
rect 49386 662458 49622 662694
rect 49706 662458 49942 662694
rect 49386 626778 49622 627014
rect 49706 626778 49942 627014
rect 49386 626458 49622 626694
rect 49706 626458 49942 626694
rect 49386 590778 49622 591014
rect 49706 590778 49942 591014
rect 49386 590458 49622 590694
rect 49706 590458 49942 590694
rect 49386 554778 49622 555014
rect 49706 554778 49942 555014
rect 49386 554458 49622 554694
rect 49706 554458 49942 554694
rect 49386 518778 49622 519014
rect 49706 518778 49942 519014
rect 49386 518458 49622 518694
rect 49706 518458 49942 518694
rect 49386 482778 49622 483014
rect 49706 482778 49942 483014
rect 49386 482458 49622 482694
rect 49706 482458 49942 482694
rect 49386 446778 49622 447014
rect 49706 446778 49942 447014
rect 49386 446458 49622 446694
rect 49706 446458 49942 446694
rect 49386 410778 49622 411014
rect 49706 410778 49942 411014
rect 49386 410458 49622 410694
rect 49706 410458 49942 410694
rect 49386 374778 49622 375014
rect 49706 374778 49942 375014
rect 49386 374458 49622 374694
rect 49706 374458 49942 374694
rect 49386 338778 49622 339014
rect 49706 338778 49942 339014
rect 49386 338458 49622 338694
rect 49706 338458 49942 338694
rect 49386 302778 49622 303014
rect 49706 302778 49942 303014
rect 49386 302458 49622 302694
rect 49706 302458 49942 302694
rect 49386 266778 49622 267014
rect 49706 266778 49942 267014
rect 49386 266458 49622 266694
rect 49706 266458 49942 266694
rect 49386 230778 49622 231014
rect 49706 230778 49942 231014
rect 49386 230458 49622 230694
rect 49706 230458 49942 230694
rect 49386 194778 49622 195014
rect 49706 194778 49942 195014
rect 49386 194458 49622 194694
rect 49706 194458 49942 194694
rect 49386 158778 49622 159014
rect 49706 158778 49942 159014
rect 49386 158458 49622 158694
rect 49706 158458 49942 158694
rect 49386 122778 49622 123014
rect 49706 122778 49942 123014
rect 49386 122458 49622 122694
rect 49706 122458 49942 122694
rect 49386 86778 49622 87014
rect 49706 86778 49942 87014
rect 49386 86458 49622 86694
rect 49706 86458 49942 86694
rect 49386 50778 49622 51014
rect 49706 50778 49942 51014
rect 49386 50458 49622 50694
rect 49706 50458 49942 50694
rect 49386 14778 49622 15014
rect 49706 14778 49942 15014
rect 49386 14458 49622 14694
rect 49706 14458 49942 14694
rect 49386 -3462 49622 -3226
rect 49706 -3462 49942 -3226
rect 49386 -3782 49622 -3546
rect 49706 -3782 49942 -3546
rect 53106 708442 53342 708678
rect 53426 708442 53662 708678
rect 53106 708122 53342 708358
rect 53426 708122 53662 708358
rect 53106 666498 53342 666734
rect 53426 666498 53662 666734
rect 53106 666178 53342 666414
rect 53426 666178 53662 666414
rect 53106 630498 53342 630734
rect 53426 630498 53662 630734
rect 53106 630178 53342 630414
rect 53426 630178 53662 630414
rect 53106 594498 53342 594734
rect 53426 594498 53662 594734
rect 53106 594178 53342 594414
rect 53426 594178 53662 594414
rect 53106 558498 53342 558734
rect 53426 558498 53662 558734
rect 53106 558178 53342 558414
rect 53426 558178 53662 558414
rect 53106 522498 53342 522734
rect 53426 522498 53662 522734
rect 53106 522178 53342 522414
rect 53426 522178 53662 522414
rect 53106 486498 53342 486734
rect 53426 486498 53662 486734
rect 53106 486178 53342 486414
rect 53426 486178 53662 486414
rect 53106 450498 53342 450734
rect 53426 450498 53662 450734
rect 53106 450178 53342 450414
rect 53426 450178 53662 450414
rect 53106 414498 53342 414734
rect 53426 414498 53662 414734
rect 53106 414178 53342 414414
rect 53426 414178 53662 414414
rect 53106 378498 53342 378734
rect 53426 378498 53662 378734
rect 53106 378178 53342 378414
rect 53426 378178 53662 378414
rect 53106 342498 53342 342734
rect 53426 342498 53662 342734
rect 53106 342178 53342 342414
rect 53426 342178 53662 342414
rect 53106 306498 53342 306734
rect 53426 306498 53662 306734
rect 53106 306178 53342 306414
rect 53426 306178 53662 306414
rect 53106 270498 53342 270734
rect 53426 270498 53662 270734
rect 53106 270178 53342 270414
rect 53426 270178 53662 270414
rect 53106 234498 53342 234734
rect 53426 234498 53662 234734
rect 53106 234178 53342 234414
rect 53426 234178 53662 234414
rect 53106 198498 53342 198734
rect 53426 198498 53662 198734
rect 53106 198178 53342 198414
rect 53426 198178 53662 198414
rect 53106 162498 53342 162734
rect 53426 162498 53662 162734
rect 53106 162178 53342 162414
rect 53426 162178 53662 162414
rect 53106 126498 53342 126734
rect 53426 126498 53662 126734
rect 53106 126178 53342 126414
rect 53426 126178 53662 126414
rect 53106 90498 53342 90734
rect 53426 90498 53662 90734
rect 53106 90178 53342 90414
rect 53426 90178 53662 90414
rect 53106 54498 53342 54734
rect 53426 54498 53662 54734
rect 53106 54178 53342 54414
rect 53426 54178 53662 54414
rect 53106 18498 53342 18734
rect 53426 18498 53662 18734
rect 53106 18178 53342 18414
rect 53426 18178 53662 18414
rect 53106 -4422 53342 -4186
rect 53426 -4422 53662 -4186
rect 53106 -4742 53342 -4506
rect 53426 -4742 53662 -4506
rect 56826 709402 57062 709638
rect 57146 709402 57382 709638
rect 56826 709082 57062 709318
rect 57146 709082 57382 709318
rect 56826 670218 57062 670454
rect 57146 670218 57382 670454
rect 56826 669898 57062 670134
rect 57146 669898 57382 670134
rect 56826 634218 57062 634454
rect 57146 634218 57382 634454
rect 56826 633898 57062 634134
rect 57146 633898 57382 634134
rect 56826 598218 57062 598454
rect 57146 598218 57382 598454
rect 56826 597898 57062 598134
rect 57146 597898 57382 598134
rect 56826 562218 57062 562454
rect 57146 562218 57382 562454
rect 56826 561898 57062 562134
rect 57146 561898 57382 562134
rect 56826 526218 57062 526454
rect 57146 526218 57382 526454
rect 56826 525898 57062 526134
rect 57146 525898 57382 526134
rect 56826 490218 57062 490454
rect 57146 490218 57382 490454
rect 56826 489898 57062 490134
rect 57146 489898 57382 490134
rect 56826 454218 57062 454454
rect 57146 454218 57382 454454
rect 56826 453898 57062 454134
rect 57146 453898 57382 454134
rect 56826 418218 57062 418454
rect 57146 418218 57382 418454
rect 56826 417898 57062 418134
rect 57146 417898 57382 418134
rect 56826 382218 57062 382454
rect 57146 382218 57382 382454
rect 56826 381898 57062 382134
rect 57146 381898 57382 382134
rect 56826 346218 57062 346454
rect 57146 346218 57382 346454
rect 56826 345898 57062 346134
rect 57146 345898 57382 346134
rect 56826 310218 57062 310454
rect 57146 310218 57382 310454
rect 56826 309898 57062 310134
rect 57146 309898 57382 310134
rect 56826 274218 57062 274454
rect 57146 274218 57382 274454
rect 56826 273898 57062 274134
rect 57146 273898 57382 274134
rect 56826 238218 57062 238454
rect 57146 238218 57382 238454
rect 56826 237898 57062 238134
rect 57146 237898 57382 238134
rect 56826 202218 57062 202454
rect 57146 202218 57382 202454
rect 56826 201898 57062 202134
rect 57146 201898 57382 202134
rect 56826 166218 57062 166454
rect 57146 166218 57382 166454
rect 56826 165898 57062 166134
rect 57146 165898 57382 166134
rect 56826 130218 57062 130454
rect 57146 130218 57382 130454
rect 56826 129898 57062 130134
rect 57146 129898 57382 130134
rect 56826 94218 57062 94454
rect 57146 94218 57382 94454
rect 56826 93898 57062 94134
rect 57146 93898 57382 94134
rect 56826 58218 57062 58454
rect 57146 58218 57382 58454
rect 56826 57898 57062 58134
rect 57146 57898 57382 58134
rect 56826 22218 57062 22454
rect 57146 22218 57382 22454
rect 56826 21898 57062 22134
rect 57146 21898 57382 22134
rect 60546 710362 60782 710598
rect 60866 710362 61102 710598
rect 60546 710042 60782 710278
rect 60866 710042 61102 710278
rect 60546 673938 60782 674174
rect 60866 673938 61102 674174
rect 60546 673618 60782 673854
rect 60866 673618 61102 673854
rect 60546 637938 60782 638174
rect 60866 637938 61102 638174
rect 60546 637618 60782 637854
rect 60866 637618 61102 637854
rect 60546 601938 60782 602174
rect 60866 601938 61102 602174
rect 60546 601618 60782 601854
rect 60866 601618 61102 601854
rect 60546 565938 60782 566174
rect 60866 565938 61102 566174
rect 60546 565618 60782 565854
rect 60866 565618 61102 565854
rect 60546 529938 60782 530174
rect 60866 529938 61102 530174
rect 60546 529618 60782 529854
rect 60866 529618 61102 529854
rect 60546 493938 60782 494174
rect 60866 493938 61102 494174
rect 60546 493618 60782 493854
rect 60866 493618 61102 493854
rect 60546 457938 60782 458174
rect 60866 457938 61102 458174
rect 60546 457618 60782 457854
rect 60866 457618 61102 457854
rect 60546 421938 60782 422174
rect 60866 421938 61102 422174
rect 60546 421618 60782 421854
rect 60866 421618 61102 421854
rect 60546 385938 60782 386174
rect 60866 385938 61102 386174
rect 60546 385618 60782 385854
rect 60866 385618 61102 385854
rect 60546 349938 60782 350174
rect 60866 349938 61102 350174
rect 60546 349618 60782 349854
rect 60866 349618 61102 349854
rect 60546 313938 60782 314174
rect 60866 313938 61102 314174
rect 60546 313618 60782 313854
rect 60866 313618 61102 313854
rect 60546 277938 60782 278174
rect 60866 277938 61102 278174
rect 60546 277618 60782 277854
rect 60866 277618 61102 277854
rect 60546 241938 60782 242174
rect 60866 241938 61102 242174
rect 60546 241618 60782 241854
rect 60866 241618 61102 241854
rect 60546 205938 60782 206174
rect 60866 205938 61102 206174
rect 60546 205618 60782 205854
rect 60866 205618 61102 205854
rect 60546 169938 60782 170174
rect 60866 169938 61102 170174
rect 60546 169618 60782 169854
rect 60866 169618 61102 169854
rect 60546 133938 60782 134174
rect 60866 133938 61102 134174
rect 60546 133618 60782 133854
rect 60866 133618 61102 133854
rect 60546 97938 60782 98174
rect 60866 97938 61102 98174
rect 60546 97618 60782 97854
rect 60866 97618 61102 97854
rect 60546 61938 60782 62174
rect 60866 61938 61102 62174
rect 60546 61618 60782 61854
rect 60866 61618 61102 61854
rect 60546 25938 60782 26174
rect 60866 25938 61102 26174
rect 60546 25618 60782 25854
rect 60866 25618 61102 25854
rect 57750 11782 57986 12018
rect 56826 -5382 57062 -5146
rect 57146 -5382 57382 -5146
rect 56826 -5702 57062 -5466
rect 57146 -5702 57382 -5466
rect 60546 -6342 60782 -6106
rect 60866 -6342 61102 -6106
rect 60546 -6662 60782 -6426
rect 60866 -6662 61102 -6426
rect 64266 711322 64502 711558
rect 64586 711322 64822 711558
rect 64266 711002 64502 711238
rect 64586 711002 64822 711238
rect 64266 677658 64502 677894
rect 64586 677658 64822 677894
rect 64266 677338 64502 677574
rect 64586 677338 64822 677574
rect 64266 641658 64502 641894
rect 64586 641658 64822 641894
rect 64266 641338 64502 641574
rect 64586 641338 64822 641574
rect 64266 605658 64502 605894
rect 64586 605658 64822 605894
rect 64266 605338 64502 605574
rect 64586 605338 64822 605574
rect 64266 569658 64502 569894
rect 64586 569658 64822 569894
rect 64266 569338 64502 569574
rect 64586 569338 64822 569574
rect 64266 533658 64502 533894
rect 64586 533658 64822 533894
rect 64266 533338 64502 533574
rect 64586 533338 64822 533574
rect 64266 497658 64502 497894
rect 64586 497658 64822 497894
rect 64266 497338 64502 497574
rect 64586 497338 64822 497574
rect 64266 461658 64502 461894
rect 64586 461658 64822 461894
rect 64266 461338 64502 461574
rect 64586 461338 64822 461574
rect 64266 425658 64502 425894
rect 64586 425658 64822 425894
rect 64266 425338 64502 425574
rect 64586 425338 64822 425574
rect 64266 389658 64502 389894
rect 64586 389658 64822 389894
rect 64266 389338 64502 389574
rect 64586 389338 64822 389574
rect 64266 353658 64502 353894
rect 64586 353658 64822 353894
rect 64266 353338 64502 353574
rect 64586 353338 64822 353574
rect 64266 317658 64502 317894
rect 64586 317658 64822 317894
rect 64266 317338 64502 317574
rect 64586 317338 64822 317574
rect 64266 281658 64502 281894
rect 64586 281658 64822 281894
rect 64266 281338 64502 281574
rect 64586 281338 64822 281574
rect 64266 245658 64502 245894
rect 64586 245658 64822 245894
rect 64266 245338 64502 245574
rect 64586 245338 64822 245574
rect 64266 209658 64502 209894
rect 64586 209658 64822 209894
rect 64266 209338 64502 209574
rect 64586 209338 64822 209574
rect 64266 173658 64502 173894
rect 64586 173658 64822 173894
rect 64266 173338 64502 173574
rect 64586 173338 64822 173574
rect 64266 137658 64502 137894
rect 64586 137658 64822 137894
rect 64266 137338 64502 137574
rect 64586 137338 64822 137574
rect 64266 101658 64502 101894
rect 64586 101658 64822 101894
rect 64266 101338 64502 101574
rect 64586 101338 64822 101574
rect 64266 65658 64502 65894
rect 64586 65658 64822 65894
rect 64266 65338 64502 65574
rect 64586 65338 64822 65574
rect 64266 29658 64502 29894
rect 64586 29658 64822 29894
rect 64266 29338 64502 29574
rect 64586 29338 64822 29574
rect 74226 704602 74462 704838
rect 74546 704602 74782 704838
rect 74226 704282 74462 704518
rect 74546 704282 74782 704518
rect 74226 687618 74462 687854
rect 74546 687618 74782 687854
rect 74226 687298 74462 687534
rect 74546 687298 74782 687534
rect 74226 651618 74462 651854
rect 74546 651618 74782 651854
rect 74226 651298 74462 651534
rect 74546 651298 74782 651534
rect 74226 615618 74462 615854
rect 74546 615618 74782 615854
rect 74226 615298 74462 615534
rect 74546 615298 74782 615534
rect 74226 579618 74462 579854
rect 74546 579618 74782 579854
rect 74226 579298 74462 579534
rect 74546 579298 74782 579534
rect 74226 543618 74462 543854
rect 74546 543618 74782 543854
rect 74226 543298 74462 543534
rect 74546 543298 74782 543534
rect 74226 507618 74462 507854
rect 74546 507618 74782 507854
rect 74226 507298 74462 507534
rect 74546 507298 74782 507534
rect 74226 471618 74462 471854
rect 74546 471618 74782 471854
rect 74226 471298 74462 471534
rect 74546 471298 74782 471534
rect 74226 435618 74462 435854
rect 74546 435618 74782 435854
rect 74226 435298 74462 435534
rect 74546 435298 74782 435534
rect 74226 399618 74462 399854
rect 74546 399618 74782 399854
rect 74226 399298 74462 399534
rect 74546 399298 74782 399534
rect 74226 363618 74462 363854
rect 74546 363618 74782 363854
rect 74226 363298 74462 363534
rect 74546 363298 74782 363534
rect 74226 327618 74462 327854
rect 74546 327618 74782 327854
rect 74226 327298 74462 327534
rect 74546 327298 74782 327534
rect 74226 291618 74462 291854
rect 74546 291618 74782 291854
rect 74226 291298 74462 291534
rect 74546 291298 74782 291534
rect 74226 255618 74462 255854
rect 74546 255618 74782 255854
rect 74226 255298 74462 255534
rect 74546 255298 74782 255534
rect 74226 219618 74462 219854
rect 74546 219618 74782 219854
rect 74226 219298 74462 219534
rect 74546 219298 74782 219534
rect 74226 183618 74462 183854
rect 74546 183618 74782 183854
rect 74226 183298 74462 183534
rect 74546 183298 74782 183534
rect 74226 147618 74462 147854
rect 74546 147618 74782 147854
rect 74226 147298 74462 147534
rect 74546 147298 74782 147534
rect 74226 111618 74462 111854
rect 74546 111618 74782 111854
rect 74226 111298 74462 111534
rect 74546 111298 74782 111534
rect 74226 75618 74462 75854
rect 74546 75618 74782 75854
rect 74226 75298 74462 75534
rect 74546 75298 74782 75534
rect 74226 39618 74462 39854
rect 74546 39618 74782 39854
rect 74226 39298 74462 39534
rect 74546 39298 74782 39534
rect 67318 8382 67554 8618
rect 77946 705562 78182 705798
rect 78266 705562 78502 705798
rect 77946 705242 78182 705478
rect 78266 705242 78502 705478
rect 77946 691338 78182 691574
rect 78266 691338 78502 691574
rect 77946 691018 78182 691254
rect 78266 691018 78502 691254
rect 77946 655338 78182 655574
rect 78266 655338 78502 655574
rect 77946 655018 78182 655254
rect 78266 655018 78502 655254
rect 77946 619338 78182 619574
rect 78266 619338 78502 619574
rect 77946 619018 78182 619254
rect 78266 619018 78502 619254
rect 77946 583338 78182 583574
rect 78266 583338 78502 583574
rect 77946 583018 78182 583254
rect 78266 583018 78502 583254
rect 77946 547338 78182 547574
rect 78266 547338 78502 547574
rect 77946 547018 78182 547254
rect 78266 547018 78502 547254
rect 77946 511338 78182 511574
rect 78266 511338 78502 511574
rect 77946 511018 78182 511254
rect 78266 511018 78502 511254
rect 77946 475338 78182 475574
rect 78266 475338 78502 475574
rect 77946 475018 78182 475254
rect 78266 475018 78502 475254
rect 77946 439338 78182 439574
rect 78266 439338 78502 439574
rect 77946 439018 78182 439254
rect 78266 439018 78502 439254
rect 77946 403338 78182 403574
rect 78266 403338 78502 403574
rect 77946 403018 78182 403254
rect 78266 403018 78502 403254
rect 77946 367338 78182 367574
rect 78266 367338 78502 367574
rect 77946 367018 78182 367254
rect 78266 367018 78502 367254
rect 77946 331338 78182 331574
rect 78266 331338 78502 331574
rect 77946 331018 78182 331254
rect 78266 331018 78502 331254
rect 77946 295338 78182 295574
rect 78266 295338 78502 295574
rect 77946 295018 78182 295254
rect 78266 295018 78502 295254
rect 77946 259338 78182 259574
rect 78266 259338 78502 259574
rect 77946 259018 78182 259254
rect 78266 259018 78502 259254
rect 77946 223338 78182 223574
rect 78266 223338 78502 223574
rect 77946 223018 78182 223254
rect 78266 223018 78502 223254
rect 77946 187338 78182 187574
rect 78266 187338 78502 187574
rect 77946 187018 78182 187254
rect 78266 187018 78502 187254
rect 77946 151338 78182 151574
rect 78266 151338 78502 151574
rect 77946 151018 78182 151254
rect 78266 151018 78502 151254
rect 77946 115338 78182 115574
rect 78266 115338 78502 115574
rect 77946 115018 78182 115254
rect 78266 115018 78502 115254
rect 77946 79338 78182 79574
rect 78266 79338 78502 79574
rect 77946 79018 78182 79254
rect 78266 79018 78502 79254
rect 77946 43338 78182 43574
rect 78266 43338 78502 43574
rect 77946 43018 78182 43254
rect 78266 43018 78502 43254
rect 77946 7338 78182 7574
rect 78266 7338 78502 7574
rect 77946 7018 78182 7254
rect 78266 7018 78502 7254
rect 74226 3618 74462 3854
rect 74546 3618 74782 3854
rect 74226 3298 74462 3534
rect 74546 3298 74782 3534
rect 64266 -7302 64502 -7066
rect 64586 -7302 64822 -7066
rect 64266 -7622 64502 -7386
rect 64586 -7622 64822 -7386
rect 74226 -582 74462 -346
rect 74546 -582 74782 -346
rect 74226 -902 74462 -666
rect 74546 -902 74782 -666
rect 77946 -1542 78182 -1306
rect 78266 -1542 78502 -1306
rect 77946 -1862 78182 -1626
rect 78266 -1862 78502 -1626
rect 81666 706522 81902 706758
rect 81986 706522 82222 706758
rect 81666 706202 81902 706438
rect 81986 706202 82222 706438
rect 81666 695058 81902 695294
rect 81986 695058 82222 695294
rect 81666 694738 81902 694974
rect 81986 694738 82222 694974
rect 81666 659058 81902 659294
rect 81986 659058 82222 659294
rect 81666 658738 81902 658974
rect 81986 658738 82222 658974
rect 81666 623058 81902 623294
rect 81986 623058 82222 623294
rect 81666 622738 81902 622974
rect 81986 622738 82222 622974
rect 81666 587058 81902 587294
rect 81986 587058 82222 587294
rect 81666 586738 81902 586974
rect 81986 586738 82222 586974
rect 81666 551058 81902 551294
rect 81986 551058 82222 551294
rect 81666 550738 81902 550974
rect 81986 550738 82222 550974
rect 81666 515058 81902 515294
rect 81986 515058 82222 515294
rect 81666 514738 81902 514974
rect 81986 514738 82222 514974
rect 81666 479058 81902 479294
rect 81986 479058 82222 479294
rect 81666 478738 81902 478974
rect 81986 478738 82222 478974
rect 81666 443058 81902 443294
rect 81986 443058 82222 443294
rect 81666 442738 81902 442974
rect 81986 442738 82222 442974
rect 81666 407058 81902 407294
rect 81986 407058 82222 407294
rect 81666 406738 81902 406974
rect 81986 406738 82222 406974
rect 81666 371058 81902 371294
rect 81986 371058 82222 371294
rect 81666 370738 81902 370974
rect 81986 370738 82222 370974
rect 81666 335058 81902 335294
rect 81986 335058 82222 335294
rect 81666 334738 81902 334974
rect 81986 334738 82222 334974
rect 81666 299058 81902 299294
rect 81986 299058 82222 299294
rect 81666 298738 81902 298974
rect 81986 298738 82222 298974
rect 81666 263058 81902 263294
rect 81986 263058 82222 263294
rect 81666 262738 81902 262974
rect 81986 262738 82222 262974
rect 81666 227058 81902 227294
rect 81986 227058 82222 227294
rect 81666 226738 81902 226974
rect 81986 226738 82222 226974
rect 81666 191058 81902 191294
rect 81986 191058 82222 191294
rect 81666 190738 81902 190974
rect 81986 190738 82222 190974
rect 85386 707482 85622 707718
rect 85706 707482 85942 707718
rect 85386 707162 85622 707398
rect 85706 707162 85942 707398
rect 85386 698778 85622 699014
rect 85706 698778 85942 699014
rect 85386 698458 85622 698694
rect 85706 698458 85942 698694
rect 85386 662778 85622 663014
rect 85706 662778 85942 663014
rect 85386 662458 85622 662694
rect 85706 662458 85942 662694
rect 85386 626778 85622 627014
rect 85706 626778 85942 627014
rect 85386 626458 85622 626694
rect 85706 626458 85942 626694
rect 85386 590778 85622 591014
rect 85706 590778 85942 591014
rect 85386 590458 85622 590694
rect 85706 590458 85942 590694
rect 85386 554778 85622 555014
rect 85706 554778 85942 555014
rect 85386 554458 85622 554694
rect 85706 554458 85942 554694
rect 85386 518778 85622 519014
rect 85706 518778 85942 519014
rect 85386 518458 85622 518694
rect 85706 518458 85942 518694
rect 85386 482778 85622 483014
rect 85706 482778 85942 483014
rect 85386 482458 85622 482694
rect 85706 482458 85942 482694
rect 85386 446778 85622 447014
rect 85706 446778 85942 447014
rect 85386 446458 85622 446694
rect 85706 446458 85942 446694
rect 85386 410778 85622 411014
rect 85706 410778 85942 411014
rect 85386 410458 85622 410694
rect 85706 410458 85942 410694
rect 85386 374778 85622 375014
rect 85706 374778 85942 375014
rect 85386 374458 85622 374694
rect 85706 374458 85942 374694
rect 85386 338778 85622 339014
rect 85706 338778 85942 339014
rect 85386 338458 85622 338694
rect 85706 338458 85942 338694
rect 85386 302778 85622 303014
rect 85706 302778 85942 303014
rect 85386 302458 85622 302694
rect 85706 302458 85942 302694
rect 85386 266778 85622 267014
rect 85706 266778 85942 267014
rect 85386 266458 85622 266694
rect 85706 266458 85942 266694
rect 85386 230778 85622 231014
rect 85706 230778 85942 231014
rect 85386 230458 85622 230694
rect 85706 230458 85942 230694
rect 85386 194778 85622 195014
rect 85706 194778 85942 195014
rect 85386 194458 85622 194694
rect 85706 194458 85942 194694
rect 84250 183618 84486 183854
rect 84250 183298 84486 183534
rect 81666 155058 81902 155294
rect 81986 155058 82222 155294
rect 81666 154738 81902 154974
rect 81986 154738 82222 154974
rect 85386 158778 85622 159014
rect 85706 158778 85942 159014
rect 85386 158458 85622 158694
rect 85706 158458 85942 158694
rect 84250 147618 84486 147854
rect 84250 147298 84486 147534
rect 81666 119058 81902 119294
rect 81986 119058 82222 119294
rect 81666 118738 81902 118974
rect 81986 118738 82222 118974
rect 85386 122778 85622 123014
rect 85706 122778 85942 123014
rect 85386 122458 85622 122694
rect 85706 122458 85942 122694
rect 84250 111618 84486 111854
rect 84250 111298 84486 111534
rect 81666 83058 81902 83294
rect 81986 83058 82222 83294
rect 81666 82738 81902 82974
rect 81986 82738 82222 82974
rect 81666 47058 81902 47294
rect 81986 47058 82222 47294
rect 81666 46738 81902 46974
rect 81986 46738 82222 46974
rect 81666 11058 81902 11294
rect 81986 11058 82222 11294
rect 81666 10738 81902 10974
rect 81986 10738 82222 10974
rect 81666 -2502 81902 -2266
rect 81986 -2502 82222 -2266
rect 81666 -2822 81902 -2586
rect 81986 -2822 82222 -2586
rect 85386 86778 85622 87014
rect 85706 86778 85942 87014
rect 85386 86458 85622 86694
rect 85706 86458 85942 86694
rect 85386 50778 85622 51014
rect 85706 50778 85942 51014
rect 85386 50458 85622 50694
rect 85706 50458 85942 50694
rect 85386 14778 85622 15014
rect 85706 14778 85942 15014
rect 85386 14458 85622 14694
rect 85706 14458 85942 14694
rect 85386 -3462 85622 -3226
rect 85706 -3462 85942 -3226
rect 85386 -3782 85622 -3546
rect 85706 -3782 85942 -3546
rect 89106 708442 89342 708678
rect 89426 708442 89662 708678
rect 89106 708122 89342 708358
rect 89426 708122 89662 708358
rect 89106 666498 89342 666734
rect 89426 666498 89662 666734
rect 89106 666178 89342 666414
rect 89426 666178 89662 666414
rect 89106 630498 89342 630734
rect 89426 630498 89662 630734
rect 89106 630178 89342 630414
rect 89426 630178 89662 630414
rect 89106 594498 89342 594734
rect 89426 594498 89662 594734
rect 89106 594178 89342 594414
rect 89426 594178 89662 594414
rect 89106 558498 89342 558734
rect 89426 558498 89662 558734
rect 89106 558178 89342 558414
rect 89426 558178 89662 558414
rect 89106 522498 89342 522734
rect 89426 522498 89662 522734
rect 89106 522178 89342 522414
rect 89426 522178 89662 522414
rect 89106 486498 89342 486734
rect 89426 486498 89662 486734
rect 89106 486178 89342 486414
rect 89426 486178 89662 486414
rect 89106 450498 89342 450734
rect 89426 450498 89662 450734
rect 89106 450178 89342 450414
rect 89426 450178 89662 450414
rect 89106 414498 89342 414734
rect 89426 414498 89662 414734
rect 89106 414178 89342 414414
rect 89426 414178 89662 414414
rect 89106 378498 89342 378734
rect 89426 378498 89662 378734
rect 89106 378178 89342 378414
rect 89426 378178 89662 378414
rect 89106 342498 89342 342734
rect 89426 342498 89662 342734
rect 89106 342178 89342 342414
rect 89426 342178 89662 342414
rect 89106 306498 89342 306734
rect 89426 306498 89662 306734
rect 89106 306178 89342 306414
rect 89426 306178 89662 306414
rect 89106 270498 89342 270734
rect 89426 270498 89662 270734
rect 89106 270178 89342 270414
rect 89426 270178 89662 270414
rect 89106 234498 89342 234734
rect 89426 234498 89662 234734
rect 89106 234178 89342 234414
rect 89426 234178 89662 234414
rect 89106 198498 89342 198734
rect 89426 198498 89662 198734
rect 89106 198178 89342 198414
rect 89426 198178 89662 198414
rect 89106 162498 89342 162734
rect 89426 162498 89662 162734
rect 89106 162178 89342 162414
rect 89426 162178 89662 162414
rect 89106 126498 89342 126734
rect 89426 126498 89662 126734
rect 89106 126178 89342 126414
rect 89426 126178 89662 126414
rect 89106 90498 89342 90734
rect 89426 90498 89662 90734
rect 89106 90178 89342 90414
rect 89426 90178 89662 90414
rect 92826 709402 93062 709638
rect 93146 709402 93382 709638
rect 92826 709082 93062 709318
rect 93146 709082 93382 709318
rect 92826 670218 93062 670454
rect 93146 670218 93382 670454
rect 92826 669898 93062 670134
rect 93146 669898 93382 670134
rect 92826 634218 93062 634454
rect 93146 634218 93382 634454
rect 92826 633898 93062 634134
rect 93146 633898 93382 634134
rect 92826 598218 93062 598454
rect 93146 598218 93382 598454
rect 92826 597898 93062 598134
rect 93146 597898 93382 598134
rect 92826 562218 93062 562454
rect 93146 562218 93382 562454
rect 92826 561898 93062 562134
rect 93146 561898 93382 562134
rect 92826 526218 93062 526454
rect 93146 526218 93382 526454
rect 92826 525898 93062 526134
rect 93146 525898 93382 526134
rect 92826 490218 93062 490454
rect 93146 490218 93382 490454
rect 92826 489898 93062 490134
rect 93146 489898 93382 490134
rect 92826 454218 93062 454454
rect 93146 454218 93382 454454
rect 92826 453898 93062 454134
rect 93146 453898 93382 454134
rect 92826 418218 93062 418454
rect 93146 418218 93382 418454
rect 92826 417898 93062 418134
rect 93146 417898 93382 418134
rect 92826 382218 93062 382454
rect 93146 382218 93382 382454
rect 92826 381898 93062 382134
rect 93146 381898 93382 382134
rect 92826 346218 93062 346454
rect 93146 346218 93382 346454
rect 92826 345898 93062 346134
rect 93146 345898 93382 346134
rect 92826 310218 93062 310454
rect 93146 310218 93382 310454
rect 92826 309898 93062 310134
rect 93146 309898 93382 310134
rect 92826 274218 93062 274454
rect 93146 274218 93382 274454
rect 92826 273898 93062 274134
rect 93146 273898 93382 274134
rect 92826 238218 93062 238454
rect 93146 238218 93382 238454
rect 92826 237898 93062 238134
rect 93146 237898 93382 238134
rect 92826 202218 93062 202454
rect 93146 202218 93382 202454
rect 92826 201898 93062 202134
rect 93146 201898 93382 202134
rect 92826 166218 93062 166454
rect 93146 166218 93382 166454
rect 92826 165898 93062 166134
rect 93146 165898 93382 166134
rect 92826 130218 93062 130454
rect 93146 130218 93382 130454
rect 92826 129898 93062 130134
rect 93146 129898 93382 130134
rect 92826 94218 93062 94454
rect 93146 94218 93382 94454
rect 92826 93898 93062 94134
rect 93146 93898 93382 94134
rect 89106 54498 89342 54734
rect 89426 54498 89662 54734
rect 89106 54178 89342 54414
rect 89426 54178 89662 54414
rect 89106 18498 89342 18734
rect 89426 18498 89662 18734
rect 89106 18178 89342 18414
rect 89426 18178 89662 18414
rect 96546 710362 96782 710598
rect 96866 710362 97102 710598
rect 96546 710042 96782 710278
rect 96866 710042 97102 710278
rect 96546 673938 96782 674174
rect 96866 673938 97102 674174
rect 96546 673618 96782 673854
rect 96866 673618 97102 673854
rect 96546 637938 96782 638174
rect 96866 637938 97102 638174
rect 96546 637618 96782 637854
rect 96866 637618 97102 637854
rect 96546 601938 96782 602174
rect 96866 601938 97102 602174
rect 96546 601618 96782 601854
rect 96866 601618 97102 601854
rect 96546 565938 96782 566174
rect 96866 565938 97102 566174
rect 96546 565618 96782 565854
rect 96866 565618 97102 565854
rect 96546 529938 96782 530174
rect 96866 529938 97102 530174
rect 96546 529618 96782 529854
rect 96866 529618 97102 529854
rect 96546 493938 96782 494174
rect 96866 493938 97102 494174
rect 96546 493618 96782 493854
rect 96866 493618 97102 493854
rect 96546 457938 96782 458174
rect 96866 457938 97102 458174
rect 96546 457618 96782 457854
rect 96866 457618 97102 457854
rect 96546 421938 96782 422174
rect 96866 421938 97102 422174
rect 96546 421618 96782 421854
rect 96866 421618 97102 421854
rect 96546 385938 96782 386174
rect 96866 385938 97102 386174
rect 96546 385618 96782 385854
rect 96866 385618 97102 385854
rect 96546 349938 96782 350174
rect 96866 349938 97102 350174
rect 96546 349618 96782 349854
rect 96866 349618 97102 349854
rect 96546 313938 96782 314174
rect 96866 313938 97102 314174
rect 96546 313618 96782 313854
rect 96866 313618 97102 313854
rect 96546 277938 96782 278174
rect 96866 277938 97102 278174
rect 96546 277618 96782 277854
rect 96866 277618 97102 277854
rect 96546 241938 96782 242174
rect 96866 241938 97102 242174
rect 96546 241618 96782 241854
rect 96866 241618 97102 241854
rect 96546 205938 96782 206174
rect 96866 205938 97102 206174
rect 96546 205618 96782 205854
rect 96866 205618 97102 205854
rect 100266 711322 100502 711558
rect 100586 711322 100822 711558
rect 100266 711002 100502 711238
rect 100586 711002 100822 711238
rect 100266 677658 100502 677894
rect 100586 677658 100822 677894
rect 100266 677338 100502 677574
rect 100586 677338 100822 677574
rect 100266 641658 100502 641894
rect 100586 641658 100822 641894
rect 100266 641338 100502 641574
rect 100586 641338 100822 641574
rect 100266 605658 100502 605894
rect 100586 605658 100822 605894
rect 100266 605338 100502 605574
rect 100586 605338 100822 605574
rect 100266 569658 100502 569894
rect 100586 569658 100822 569894
rect 100266 569338 100502 569574
rect 100586 569338 100822 569574
rect 100266 533658 100502 533894
rect 100586 533658 100822 533894
rect 100266 533338 100502 533574
rect 100586 533338 100822 533574
rect 100266 497658 100502 497894
rect 100586 497658 100822 497894
rect 100266 497338 100502 497574
rect 100586 497338 100822 497574
rect 100266 461658 100502 461894
rect 100586 461658 100822 461894
rect 100266 461338 100502 461574
rect 100586 461338 100822 461574
rect 100266 425658 100502 425894
rect 100586 425658 100822 425894
rect 100266 425338 100502 425574
rect 100586 425338 100822 425574
rect 100266 389658 100502 389894
rect 100586 389658 100822 389894
rect 100266 389338 100502 389574
rect 100586 389338 100822 389574
rect 100266 353658 100502 353894
rect 100586 353658 100822 353894
rect 100266 353338 100502 353574
rect 100586 353338 100822 353574
rect 100266 317658 100502 317894
rect 100586 317658 100822 317894
rect 100266 317338 100502 317574
rect 100586 317338 100822 317574
rect 100266 281658 100502 281894
rect 100586 281658 100822 281894
rect 100266 281338 100502 281574
rect 100586 281338 100822 281574
rect 100266 245658 100502 245894
rect 100586 245658 100822 245894
rect 100266 245338 100502 245574
rect 100586 245338 100822 245574
rect 100266 209658 100502 209894
rect 100586 209658 100822 209894
rect 100266 209338 100502 209574
rect 100586 209338 100822 209574
rect 110226 704602 110462 704838
rect 110546 704602 110782 704838
rect 110226 704282 110462 704518
rect 110546 704282 110782 704518
rect 110226 687618 110462 687854
rect 110546 687618 110782 687854
rect 110226 687298 110462 687534
rect 110546 687298 110782 687534
rect 110226 651618 110462 651854
rect 110546 651618 110782 651854
rect 110226 651298 110462 651534
rect 110546 651298 110782 651534
rect 110226 615618 110462 615854
rect 110546 615618 110782 615854
rect 110226 615298 110462 615534
rect 110546 615298 110782 615534
rect 110226 579618 110462 579854
rect 110546 579618 110782 579854
rect 110226 579298 110462 579534
rect 110546 579298 110782 579534
rect 110226 543618 110462 543854
rect 110546 543618 110782 543854
rect 110226 543298 110462 543534
rect 110546 543298 110782 543534
rect 110226 507618 110462 507854
rect 110546 507618 110782 507854
rect 110226 507298 110462 507534
rect 110546 507298 110782 507534
rect 110226 471618 110462 471854
rect 110546 471618 110782 471854
rect 110226 471298 110462 471534
rect 110546 471298 110782 471534
rect 110226 435618 110462 435854
rect 110546 435618 110782 435854
rect 110226 435298 110462 435534
rect 110546 435298 110782 435534
rect 110226 399618 110462 399854
rect 110546 399618 110782 399854
rect 110226 399298 110462 399534
rect 110546 399298 110782 399534
rect 110226 363618 110462 363854
rect 110546 363618 110782 363854
rect 110226 363298 110462 363534
rect 110546 363298 110782 363534
rect 110226 327618 110462 327854
rect 110546 327618 110782 327854
rect 110226 327298 110462 327534
rect 110546 327298 110782 327534
rect 110226 291618 110462 291854
rect 110546 291618 110782 291854
rect 110226 291298 110462 291534
rect 110546 291298 110782 291534
rect 110226 255618 110462 255854
rect 110546 255618 110782 255854
rect 110226 255298 110462 255534
rect 110546 255298 110782 255534
rect 110226 219618 110462 219854
rect 110546 219618 110782 219854
rect 110226 219298 110462 219534
rect 110546 219298 110782 219534
rect 113946 705562 114182 705798
rect 114266 705562 114502 705798
rect 113946 705242 114182 705478
rect 114266 705242 114502 705478
rect 113946 691338 114182 691574
rect 114266 691338 114502 691574
rect 113946 691018 114182 691254
rect 114266 691018 114502 691254
rect 113946 655338 114182 655574
rect 114266 655338 114502 655574
rect 113946 655018 114182 655254
rect 114266 655018 114502 655254
rect 113946 619338 114182 619574
rect 114266 619338 114502 619574
rect 113946 619018 114182 619254
rect 114266 619018 114502 619254
rect 113946 583338 114182 583574
rect 114266 583338 114502 583574
rect 113946 583018 114182 583254
rect 114266 583018 114502 583254
rect 113946 547338 114182 547574
rect 114266 547338 114502 547574
rect 113946 547018 114182 547254
rect 114266 547018 114502 547254
rect 113946 511338 114182 511574
rect 114266 511338 114502 511574
rect 113946 511018 114182 511254
rect 114266 511018 114502 511254
rect 113946 475338 114182 475574
rect 114266 475338 114502 475574
rect 113946 475018 114182 475254
rect 114266 475018 114502 475254
rect 113946 439338 114182 439574
rect 114266 439338 114502 439574
rect 113946 439018 114182 439254
rect 114266 439018 114502 439254
rect 113946 403338 114182 403574
rect 114266 403338 114502 403574
rect 113946 403018 114182 403254
rect 114266 403018 114502 403254
rect 113946 367338 114182 367574
rect 114266 367338 114502 367574
rect 113946 367018 114182 367254
rect 114266 367018 114502 367254
rect 113946 331338 114182 331574
rect 114266 331338 114502 331574
rect 113946 331018 114182 331254
rect 114266 331018 114502 331254
rect 113946 295338 114182 295574
rect 114266 295338 114502 295574
rect 113946 295018 114182 295254
rect 114266 295018 114502 295254
rect 113946 259338 114182 259574
rect 114266 259338 114502 259574
rect 113946 259018 114182 259254
rect 114266 259018 114502 259254
rect 113946 223338 114182 223574
rect 114266 223338 114502 223574
rect 113946 223018 114182 223254
rect 114266 223018 114502 223254
rect 117666 706522 117902 706758
rect 117986 706522 118222 706758
rect 117666 706202 117902 706438
rect 117986 706202 118222 706438
rect 117666 695058 117902 695294
rect 117986 695058 118222 695294
rect 117666 694738 117902 694974
rect 117986 694738 118222 694974
rect 117666 659058 117902 659294
rect 117986 659058 118222 659294
rect 117666 658738 117902 658974
rect 117986 658738 118222 658974
rect 117666 623058 117902 623294
rect 117986 623058 118222 623294
rect 117666 622738 117902 622974
rect 117986 622738 118222 622974
rect 117666 587058 117902 587294
rect 117986 587058 118222 587294
rect 117666 586738 117902 586974
rect 117986 586738 118222 586974
rect 117666 551058 117902 551294
rect 117986 551058 118222 551294
rect 117666 550738 117902 550974
rect 117986 550738 118222 550974
rect 117666 515058 117902 515294
rect 117986 515058 118222 515294
rect 117666 514738 117902 514974
rect 117986 514738 118222 514974
rect 117666 479058 117902 479294
rect 117986 479058 118222 479294
rect 117666 478738 117902 478974
rect 117986 478738 118222 478974
rect 117666 443058 117902 443294
rect 117986 443058 118222 443294
rect 117666 442738 117902 442974
rect 117986 442738 118222 442974
rect 117666 407058 117902 407294
rect 117986 407058 118222 407294
rect 117666 406738 117902 406974
rect 117986 406738 118222 406974
rect 117666 371058 117902 371294
rect 117986 371058 118222 371294
rect 117666 370738 117902 370974
rect 117986 370738 118222 370974
rect 117666 335058 117902 335294
rect 117986 335058 118222 335294
rect 117666 334738 117902 334974
rect 117986 334738 118222 334974
rect 117666 299058 117902 299294
rect 117986 299058 118222 299294
rect 117666 298738 117902 298974
rect 117986 298738 118222 298974
rect 117666 263058 117902 263294
rect 117986 263058 118222 263294
rect 117666 262738 117902 262974
rect 117986 262738 118222 262974
rect 117666 227058 117902 227294
rect 117986 227058 118222 227294
rect 117666 226738 117902 226974
rect 117986 226738 118222 226974
rect 117666 191058 117902 191294
rect 117986 191058 118222 191294
rect 117666 190738 117902 190974
rect 117986 190738 118222 190974
rect 121386 707482 121622 707718
rect 121706 707482 121942 707718
rect 121386 707162 121622 707398
rect 121706 707162 121942 707398
rect 121386 698778 121622 699014
rect 121706 698778 121942 699014
rect 121386 698458 121622 698694
rect 121706 698458 121942 698694
rect 121386 662778 121622 663014
rect 121706 662778 121942 663014
rect 121386 662458 121622 662694
rect 121706 662458 121942 662694
rect 121386 626778 121622 627014
rect 121706 626778 121942 627014
rect 121386 626458 121622 626694
rect 121706 626458 121942 626694
rect 121386 590778 121622 591014
rect 121706 590778 121942 591014
rect 121386 590458 121622 590694
rect 121706 590458 121942 590694
rect 121386 554778 121622 555014
rect 121706 554778 121942 555014
rect 121386 554458 121622 554694
rect 121706 554458 121942 554694
rect 121386 518778 121622 519014
rect 121706 518778 121942 519014
rect 121386 518458 121622 518694
rect 121706 518458 121942 518694
rect 121386 482778 121622 483014
rect 121706 482778 121942 483014
rect 121386 482458 121622 482694
rect 121706 482458 121942 482694
rect 121386 446778 121622 447014
rect 121706 446778 121942 447014
rect 121386 446458 121622 446694
rect 121706 446458 121942 446694
rect 121386 410778 121622 411014
rect 121706 410778 121942 411014
rect 121386 410458 121622 410694
rect 121706 410458 121942 410694
rect 121386 374778 121622 375014
rect 121706 374778 121942 375014
rect 121386 374458 121622 374694
rect 121706 374458 121942 374694
rect 121386 338778 121622 339014
rect 121706 338778 121942 339014
rect 121386 338458 121622 338694
rect 121706 338458 121942 338694
rect 121386 302778 121622 303014
rect 121706 302778 121942 303014
rect 121386 302458 121622 302694
rect 121706 302458 121942 302694
rect 121386 266778 121622 267014
rect 121706 266778 121942 267014
rect 121386 266458 121622 266694
rect 121706 266458 121942 266694
rect 121386 230778 121622 231014
rect 121706 230778 121942 231014
rect 121386 230458 121622 230694
rect 121706 230458 121942 230694
rect 121386 194778 121622 195014
rect 121706 194778 121942 195014
rect 121386 194458 121622 194694
rect 121706 194458 121942 194694
rect 125106 708442 125342 708678
rect 125426 708442 125662 708678
rect 125106 708122 125342 708358
rect 125426 708122 125662 708358
rect 125106 666498 125342 666734
rect 125426 666498 125662 666734
rect 125106 666178 125342 666414
rect 125426 666178 125662 666414
rect 125106 630498 125342 630734
rect 125426 630498 125662 630734
rect 125106 630178 125342 630414
rect 125426 630178 125662 630414
rect 125106 594498 125342 594734
rect 125426 594498 125662 594734
rect 125106 594178 125342 594414
rect 125426 594178 125662 594414
rect 125106 558498 125342 558734
rect 125426 558498 125662 558734
rect 125106 558178 125342 558414
rect 125426 558178 125662 558414
rect 125106 522498 125342 522734
rect 125426 522498 125662 522734
rect 125106 522178 125342 522414
rect 125426 522178 125662 522414
rect 125106 486498 125342 486734
rect 125426 486498 125662 486734
rect 125106 486178 125342 486414
rect 125426 486178 125662 486414
rect 125106 450498 125342 450734
rect 125426 450498 125662 450734
rect 125106 450178 125342 450414
rect 125426 450178 125662 450414
rect 125106 414498 125342 414734
rect 125426 414498 125662 414734
rect 125106 414178 125342 414414
rect 125426 414178 125662 414414
rect 125106 378498 125342 378734
rect 125426 378498 125662 378734
rect 125106 378178 125342 378414
rect 125426 378178 125662 378414
rect 125106 342498 125342 342734
rect 125426 342498 125662 342734
rect 125106 342178 125342 342414
rect 125426 342178 125662 342414
rect 125106 306498 125342 306734
rect 125426 306498 125662 306734
rect 125106 306178 125342 306414
rect 125426 306178 125662 306414
rect 125106 270498 125342 270734
rect 125426 270498 125662 270734
rect 125106 270178 125342 270414
rect 125426 270178 125662 270414
rect 125106 234498 125342 234734
rect 125426 234498 125662 234734
rect 125106 234178 125342 234414
rect 125426 234178 125662 234414
rect 125106 198498 125342 198734
rect 125426 198498 125662 198734
rect 125106 198178 125342 198414
rect 125426 198178 125662 198414
rect 128826 709402 129062 709638
rect 129146 709402 129382 709638
rect 128826 709082 129062 709318
rect 129146 709082 129382 709318
rect 128826 670218 129062 670454
rect 129146 670218 129382 670454
rect 128826 669898 129062 670134
rect 129146 669898 129382 670134
rect 128826 634218 129062 634454
rect 129146 634218 129382 634454
rect 128826 633898 129062 634134
rect 129146 633898 129382 634134
rect 128826 598218 129062 598454
rect 129146 598218 129382 598454
rect 128826 597898 129062 598134
rect 129146 597898 129382 598134
rect 128826 562218 129062 562454
rect 129146 562218 129382 562454
rect 128826 561898 129062 562134
rect 129146 561898 129382 562134
rect 128826 526218 129062 526454
rect 129146 526218 129382 526454
rect 128826 525898 129062 526134
rect 129146 525898 129382 526134
rect 128826 490218 129062 490454
rect 129146 490218 129382 490454
rect 128826 489898 129062 490134
rect 129146 489898 129382 490134
rect 128826 454218 129062 454454
rect 129146 454218 129382 454454
rect 128826 453898 129062 454134
rect 129146 453898 129382 454134
rect 128826 418218 129062 418454
rect 129146 418218 129382 418454
rect 128826 417898 129062 418134
rect 129146 417898 129382 418134
rect 128826 382218 129062 382454
rect 129146 382218 129382 382454
rect 128826 381898 129062 382134
rect 129146 381898 129382 382134
rect 128826 346218 129062 346454
rect 129146 346218 129382 346454
rect 128826 345898 129062 346134
rect 129146 345898 129382 346134
rect 128826 310218 129062 310454
rect 129146 310218 129382 310454
rect 128826 309898 129062 310134
rect 129146 309898 129382 310134
rect 128826 274218 129062 274454
rect 129146 274218 129382 274454
rect 128826 273898 129062 274134
rect 129146 273898 129382 274134
rect 128826 238218 129062 238454
rect 129146 238218 129382 238454
rect 128826 237898 129062 238134
rect 129146 237898 129382 238134
rect 128826 202218 129062 202454
rect 129146 202218 129382 202454
rect 128826 201898 129062 202134
rect 129146 201898 129382 202134
rect 132546 710362 132782 710598
rect 132866 710362 133102 710598
rect 132546 710042 132782 710278
rect 132866 710042 133102 710278
rect 132546 673938 132782 674174
rect 132866 673938 133102 674174
rect 132546 673618 132782 673854
rect 132866 673618 133102 673854
rect 132546 637938 132782 638174
rect 132866 637938 133102 638174
rect 132546 637618 132782 637854
rect 132866 637618 133102 637854
rect 132546 601938 132782 602174
rect 132866 601938 133102 602174
rect 132546 601618 132782 601854
rect 132866 601618 133102 601854
rect 132546 565938 132782 566174
rect 132866 565938 133102 566174
rect 132546 565618 132782 565854
rect 132866 565618 133102 565854
rect 132546 529938 132782 530174
rect 132866 529938 133102 530174
rect 132546 529618 132782 529854
rect 132866 529618 133102 529854
rect 132546 493938 132782 494174
rect 132866 493938 133102 494174
rect 132546 493618 132782 493854
rect 132866 493618 133102 493854
rect 132546 457938 132782 458174
rect 132866 457938 133102 458174
rect 132546 457618 132782 457854
rect 132866 457618 133102 457854
rect 132546 421938 132782 422174
rect 132866 421938 133102 422174
rect 132546 421618 132782 421854
rect 132866 421618 133102 421854
rect 132546 385938 132782 386174
rect 132866 385938 133102 386174
rect 132546 385618 132782 385854
rect 132866 385618 133102 385854
rect 132546 349938 132782 350174
rect 132866 349938 133102 350174
rect 132546 349618 132782 349854
rect 132866 349618 133102 349854
rect 132546 313938 132782 314174
rect 132866 313938 133102 314174
rect 132546 313618 132782 313854
rect 132866 313618 133102 313854
rect 132546 277938 132782 278174
rect 132866 277938 133102 278174
rect 132546 277618 132782 277854
rect 132866 277618 133102 277854
rect 132546 241938 132782 242174
rect 132866 241938 133102 242174
rect 132546 241618 132782 241854
rect 132866 241618 133102 241854
rect 132546 205938 132782 206174
rect 132866 205938 133102 206174
rect 132546 205618 132782 205854
rect 132866 205618 133102 205854
rect 136266 711322 136502 711558
rect 136586 711322 136822 711558
rect 136266 711002 136502 711238
rect 136586 711002 136822 711238
rect 136266 677658 136502 677894
rect 136586 677658 136822 677894
rect 136266 677338 136502 677574
rect 136586 677338 136822 677574
rect 136266 641658 136502 641894
rect 136586 641658 136822 641894
rect 136266 641338 136502 641574
rect 136586 641338 136822 641574
rect 136266 605658 136502 605894
rect 136586 605658 136822 605894
rect 136266 605338 136502 605574
rect 136586 605338 136822 605574
rect 136266 569658 136502 569894
rect 136586 569658 136822 569894
rect 136266 569338 136502 569574
rect 136586 569338 136822 569574
rect 136266 533658 136502 533894
rect 136586 533658 136822 533894
rect 136266 533338 136502 533574
rect 136586 533338 136822 533574
rect 136266 497658 136502 497894
rect 136586 497658 136822 497894
rect 136266 497338 136502 497574
rect 136586 497338 136822 497574
rect 136266 461658 136502 461894
rect 136586 461658 136822 461894
rect 136266 461338 136502 461574
rect 136586 461338 136822 461574
rect 136266 425658 136502 425894
rect 136586 425658 136822 425894
rect 136266 425338 136502 425574
rect 136586 425338 136822 425574
rect 136266 389658 136502 389894
rect 136586 389658 136822 389894
rect 136266 389338 136502 389574
rect 136586 389338 136822 389574
rect 136266 353658 136502 353894
rect 136586 353658 136822 353894
rect 136266 353338 136502 353574
rect 136586 353338 136822 353574
rect 136266 317658 136502 317894
rect 136586 317658 136822 317894
rect 136266 317338 136502 317574
rect 136586 317338 136822 317574
rect 136266 281658 136502 281894
rect 136586 281658 136822 281894
rect 136266 281338 136502 281574
rect 136586 281338 136822 281574
rect 136266 245658 136502 245894
rect 136586 245658 136822 245894
rect 136266 245338 136502 245574
rect 136586 245338 136822 245574
rect 136266 209658 136502 209894
rect 136586 209658 136822 209894
rect 136266 209338 136502 209574
rect 136586 209338 136822 209574
rect 146226 704602 146462 704838
rect 146546 704602 146782 704838
rect 146226 704282 146462 704518
rect 146546 704282 146782 704518
rect 146226 687618 146462 687854
rect 146546 687618 146782 687854
rect 146226 687298 146462 687534
rect 146546 687298 146782 687534
rect 146226 651618 146462 651854
rect 146546 651618 146782 651854
rect 146226 651298 146462 651534
rect 146546 651298 146782 651534
rect 146226 615618 146462 615854
rect 146546 615618 146782 615854
rect 146226 615298 146462 615534
rect 146546 615298 146782 615534
rect 146226 579618 146462 579854
rect 146546 579618 146782 579854
rect 146226 579298 146462 579534
rect 146546 579298 146782 579534
rect 146226 543618 146462 543854
rect 146546 543618 146782 543854
rect 146226 543298 146462 543534
rect 146546 543298 146782 543534
rect 146226 507618 146462 507854
rect 146546 507618 146782 507854
rect 146226 507298 146462 507534
rect 146546 507298 146782 507534
rect 146226 471618 146462 471854
rect 146546 471618 146782 471854
rect 146226 471298 146462 471534
rect 146546 471298 146782 471534
rect 146226 435618 146462 435854
rect 146546 435618 146782 435854
rect 146226 435298 146462 435534
rect 146546 435298 146782 435534
rect 146226 399618 146462 399854
rect 146546 399618 146782 399854
rect 146226 399298 146462 399534
rect 146546 399298 146782 399534
rect 146226 363618 146462 363854
rect 146546 363618 146782 363854
rect 146226 363298 146462 363534
rect 146546 363298 146782 363534
rect 146226 327618 146462 327854
rect 146546 327618 146782 327854
rect 146226 327298 146462 327534
rect 146546 327298 146782 327534
rect 146226 291618 146462 291854
rect 146546 291618 146782 291854
rect 146226 291298 146462 291534
rect 146546 291298 146782 291534
rect 146226 255618 146462 255854
rect 146546 255618 146782 255854
rect 146226 255298 146462 255534
rect 146546 255298 146782 255534
rect 146226 219618 146462 219854
rect 146546 219618 146782 219854
rect 146226 219298 146462 219534
rect 146546 219298 146782 219534
rect 149946 705562 150182 705798
rect 150266 705562 150502 705798
rect 149946 705242 150182 705478
rect 150266 705242 150502 705478
rect 149946 691338 150182 691574
rect 150266 691338 150502 691574
rect 149946 691018 150182 691254
rect 150266 691018 150502 691254
rect 149946 655338 150182 655574
rect 150266 655338 150502 655574
rect 149946 655018 150182 655254
rect 150266 655018 150502 655254
rect 149946 619338 150182 619574
rect 150266 619338 150502 619574
rect 149946 619018 150182 619254
rect 150266 619018 150502 619254
rect 149946 583338 150182 583574
rect 150266 583338 150502 583574
rect 149946 583018 150182 583254
rect 150266 583018 150502 583254
rect 149946 547338 150182 547574
rect 150266 547338 150502 547574
rect 149946 547018 150182 547254
rect 150266 547018 150502 547254
rect 149946 511338 150182 511574
rect 150266 511338 150502 511574
rect 149946 511018 150182 511254
rect 150266 511018 150502 511254
rect 149946 475338 150182 475574
rect 150266 475338 150502 475574
rect 149946 475018 150182 475254
rect 150266 475018 150502 475254
rect 149946 439338 150182 439574
rect 150266 439338 150502 439574
rect 149946 439018 150182 439254
rect 150266 439018 150502 439254
rect 149946 403338 150182 403574
rect 150266 403338 150502 403574
rect 149946 403018 150182 403254
rect 150266 403018 150502 403254
rect 149946 367338 150182 367574
rect 150266 367338 150502 367574
rect 149946 367018 150182 367254
rect 150266 367018 150502 367254
rect 149946 331338 150182 331574
rect 150266 331338 150502 331574
rect 149946 331018 150182 331254
rect 150266 331018 150502 331254
rect 149946 295338 150182 295574
rect 150266 295338 150502 295574
rect 149946 295018 150182 295254
rect 150266 295018 150502 295254
rect 149946 259338 150182 259574
rect 150266 259338 150502 259574
rect 149946 259018 150182 259254
rect 150266 259018 150502 259254
rect 149946 223338 150182 223574
rect 150266 223338 150502 223574
rect 149946 223018 150182 223254
rect 150266 223018 150502 223254
rect 153666 706522 153902 706758
rect 153986 706522 154222 706758
rect 153666 706202 153902 706438
rect 153986 706202 154222 706438
rect 153666 695058 153902 695294
rect 153986 695058 154222 695294
rect 153666 694738 153902 694974
rect 153986 694738 154222 694974
rect 153666 659058 153902 659294
rect 153986 659058 154222 659294
rect 153666 658738 153902 658974
rect 153986 658738 154222 658974
rect 153666 623058 153902 623294
rect 153986 623058 154222 623294
rect 153666 622738 153902 622974
rect 153986 622738 154222 622974
rect 153666 587058 153902 587294
rect 153986 587058 154222 587294
rect 153666 586738 153902 586974
rect 153986 586738 154222 586974
rect 153666 551058 153902 551294
rect 153986 551058 154222 551294
rect 153666 550738 153902 550974
rect 153986 550738 154222 550974
rect 153666 515058 153902 515294
rect 153986 515058 154222 515294
rect 153666 514738 153902 514974
rect 153986 514738 154222 514974
rect 153666 479058 153902 479294
rect 153986 479058 154222 479294
rect 153666 478738 153902 478974
rect 153986 478738 154222 478974
rect 153666 443058 153902 443294
rect 153986 443058 154222 443294
rect 153666 442738 153902 442974
rect 153986 442738 154222 442974
rect 153666 407058 153902 407294
rect 153986 407058 154222 407294
rect 153666 406738 153902 406974
rect 153986 406738 154222 406974
rect 153666 371058 153902 371294
rect 153986 371058 154222 371294
rect 153666 370738 153902 370974
rect 153986 370738 154222 370974
rect 153666 335058 153902 335294
rect 153986 335058 154222 335294
rect 153666 334738 153902 334974
rect 153986 334738 154222 334974
rect 153666 299058 153902 299294
rect 153986 299058 154222 299294
rect 153666 298738 153902 298974
rect 153986 298738 154222 298974
rect 153666 263058 153902 263294
rect 153986 263058 154222 263294
rect 153666 262738 153902 262974
rect 153986 262738 154222 262974
rect 153666 227058 153902 227294
rect 153986 227058 154222 227294
rect 153666 226738 153902 226974
rect 153986 226738 154222 226974
rect 153666 191058 153902 191294
rect 153986 191058 154222 191294
rect 153666 190738 153902 190974
rect 153986 190738 154222 190974
rect 157386 707482 157622 707718
rect 157706 707482 157942 707718
rect 157386 707162 157622 707398
rect 157706 707162 157942 707398
rect 157386 698778 157622 699014
rect 157706 698778 157942 699014
rect 157386 698458 157622 698694
rect 157706 698458 157942 698694
rect 157386 662778 157622 663014
rect 157706 662778 157942 663014
rect 157386 662458 157622 662694
rect 157706 662458 157942 662694
rect 157386 626778 157622 627014
rect 157706 626778 157942 627014
rect 157386 626458 157622 626694
rect 157706 626458 157942 626694
rect 157386 590778 157622 591014
rect 157706 590778 157942 591014
rect 157386 590458 157622 590694
rect 157706 590458 157942 590694
rect 157386 554778 157622 555014
rect 157706 554778 157942 555014
rect 157386 554458 157622 554694
rect 157706 554458 157942 554694
rect 157386 518778 157622 519014
rect 157706 518778 157942 519014
rect 157386 518458 157622 518694
rect 157706 518458 157942 518694
rect 157386 482778 157622 483014
rect 157706 482778 157942 483014
rect 157386 482458 157622 482694
rect 157706 482458 157942 482694
rect 157386 446778 157622 447014
rect 157706 446778 157942 447014
rect 157386 446458 157622 446694
rect 157706 446458 157942 446694
rect 157386 410778 157622 411014
rect 157706 410778 157942 411014
rect 157386 410458 157622 410694
rect 157706 410458 157942 410694
rect 157386 374778 157622 375014
rect 157706 374778 157942 375014
rect 157386 374458 157622 374694
rect 157706 374458 157942 374694
rect 157386 338778 157622 339014
rect 157706 338778 157942 339014
rect 157386 338458 157622 338694
rect 157706 338458 157942 338694
rect 157386 302778 157622 303014
rect 157706 302778 157942 303014
rect 157386 302458 157622 302694
rect 157706 302458 157942 302694
rect 157386 266778 157622 267014
rect 157706 266778 157942 267014
rect 157386 266458 157622 266694
rect 157706 266458 157942 266694
rect 157386 230778 157622 231014
rect 157706 230778 157942 231014
rect 157386 230458 157622 230694
rect 157706 230458 157942 230694
rect 157386 194778 157622 195014
rect 157706 194778 157942 195014
rect 157386 194458 157622 194694
rect 157706 194458 157942 194694
rect 161106 708442 161342 708678
rect 161426 708442 161662 708678
rect 161106 708122 161342 708358
rect 161426 708122 161662 708358
rect 161106 666498 161342 666734
rect 161426 666498 161662 666734
rect 161106 666178 161342 666414
rect 161426 666178 161662 666414
rect 161106 630498 161342 630734
rect 161426 630498 161662 630734
rect 161106 630178 161342 630414
rect 161426 630178 161662 630414
rect 161106 594498 161342 594734
rect 161426 594498 161662 594734
rect 161106 594178 161342 594414
rect 161426 594178 161662 594414
rect 161106 558498 161342 558734
rect 161426 558498 161662 558734
rect 161106 558178 161342 558414
rect 161426 558178 161662 558414
rect 161106 522498 161342 522734
rect 161426 522498 161662 522734
rect 161106 522178 161342 522414
rect 161426 522178 161662 522414
rect 161106 486498 161342 486734
rect 161426 486498 161662 486734
rect 161106 486178 161342 486414
rect 161426 486178 161662 486414
rect 161106 450498 161342 450734
rect 161426 450498 161662 450734
rect 161106 450178 161342 450414
rect 161426 450178 161662 450414
rect 161106 414498 161342 414734
rect 161426 414498 161662 414734
rect 161106 414178 161342 414414
rect 161426 414178 161662 414414
rect 161106 378498 161342 378734
rect 161426 378498 161662 378734
rect 161106 378178 161342 378414
rect 161426 378178 161662 378414
rect 161106 342498 161342 342734
rect 161426 342498 161662 342734
rect 161106 342178 161342 342414
rect 161426 342178 161662 342414
rect 161106 306498 161342 306734
rect 161426 306498 161662 306734
rect 161106 306178 161342 306414
rect 161426 306178 161662 306414
rect 161106 270498 161342 270734
rect 161426 270498 161662 270734
rect 161106 270178 161342 270414
rect 161426 270178 161662 270414
rect 161106 234498 161342 234734
rect 161426 234498 161662 234734
rect 161106 234178 161342 234414
rect 161426 234178 161662 234414
rect 161106 198498 161342 198734
rect 161426 198498 161662 198734
rect 161106 198178 161342 198414
rect 161426 198178 161662 198414
rect 164826 709402 165062 709638
rect 165146 709402 165382 709638
rect 164826 709082 165062 709318
rect 165146 709082 165382 709318
rect 164826 670218 165062 670454
rect 165146 670218 165382 670454
rect 164826 669898 165062 670134
rect 165146 669898 165382 670134
rect 164826 634218 165062 634454
rect 165146 634218 165382 634454
rect 164826 633898 165062 634134
rect 165146 633898 165382 634134
rect 164826 598218 165062 598454
rect 165146 598218 165382 598454
rect 164826 597898 165062 598134
rect 165146 597898 165382 598134
rect 164826 562218 165062 562454
rect 165146 562218 165382 562454
rect 164826 561898 165062 562134
rect 165146 561898 165382 562134
rect 164826 526218 165062 526454
rect 165146 526218 165382 526454
rect 164826 525898 165062 526134
rect 165146 525898 165382 526134
rect 164826 490218 165062 490454
rect 165146 490218 165382 490454
rect 164826 489898 165062 490134
rect 165146 489898 165382 490134
rect 164826 454218 165062 454454
rect 165146 454218 165382 454454
rect 164826 453898 165062 454134
rect 165146 453898 165382 454134
rect 164826 418218 165062 418454
rect 165146 418218 165382 418454
rect 164826 417898 165062 418134
rect 165146 417898 165382 418134
rect 164826 382218 165062 382454
rect 165146 382218 165382 382454
rect 164826 381898 165062 382134
rect 165146 381898 165382 382134
rect 164826 346218 165062 346454
rect 165146 346218 165382 346454
rect 164826 345898 165062 346134
rect 165146 345898 165382 346134
rect 164826 310218 165062 310454
rect 165146 310218 165382 310454
rect 164826 309898 165062 310134
rect 165146 309898 165382 310134
rect 164826 274218 165062 274454
rect 165146 274218 165382 274454
rect 164826 273898 165062 274134
rect 165146 273898 165382 274134
rect 164826 238218 165062 238454
rect 165146 238218 165382 238454
rect 164826 237898 165062 238134
rect 165146 237898 165382 238134
rect 164826 202218 165062 202454
rect 165146 202218 165382 202454
rect 164826 201898 165062 202134
rect 165146 201898 165382 202134
rect 168546 710362 168782 710598
rect 168866 710362 169102 710598
rect 168546 710042 168782 710278
rect 168866 710042 169102 710278
rect 168546 673938 168782 674174
rect 168866 673938 169102 674174
rect 168546 673618 168782 673854
rect 168866 673618 169102 673854
rect 168546 637938 168782 638174
rect 168866 637938 169102 638174
rect 168546 637618 168782 637854
rect 168866 637618 169102 637854
rect 168546 601938 168782 602174
rect 168866 601938 169102 602174
rect 168546 601618 168782 601854
rect 168866 601618 169102 601854
rect 168546 565938 168782 566174
rect 168866 565938 169102 566174
rect 168546 565618 168782 565854
rect 168866 565618 169102 565854
rect 168546 529938 168782 530174
rect 168866 529938 169102 530174
rect 168546 529618 168782 529854
rect 168866 529618 169102 529854
rect 168546 493938 168782 494174
rect 168866 493938 169102 494174
rect 168546 493618 168782 493854
rect 168866 493618 169102 493854
rect 168546 457938 168782 458174
rect 168866 457938 169102 458174
rect 168546 457618 168782 457854
rect 168866 457618 169102 457854
rect 168546 421938 168782 422174
rect 168866 421938 169102 422174
rect 168546 421618 168782 421854
rect 168866 421618 169102 421854
rect 168546 385938 168782 386174
rect 168866 385938 169102 386174
rect 168546 385618 168782 385854
rect 168866 385618 169102 385854
rect 168546 349938 168782 350174
rect 168866 349938 169102 350174
rect 168546 349618 168782 349854
rect 168866 349618 169102 349854
rect 168546 313938 168782 314174
rect 168866 313938 169102 314174
rect 168546 313618 168782 313854
rect 168866 313618 169102 313854
rect 168546 277938 168782 278174
rect 168866 277938 169102 278174
rect 168546 277618 168782 277854
rect 168866 277618 169102 277854
rect 168546 241938 168782 242174
rect 168866 241938 169102 242174
rect 168546 241618 168782 241854
rect 168866 241618 169102 241854
rect 168546 205938 168782 206174
rect 168866 205938 169102 206174
rect 168546 205618 168782 205854
rect 168866 205618 169102 205854
rect 172266 711322 172502 711558
rect 172586 711322 172822 711558
rect 172266 711002 172502 711238
rect 172586 711002 172822 711238
rect 172266 677658 172502 677894
rect 172586 677658 172822 677894
rect 172266 677338 172502 677574
rect 172586 677338 172822 677574
rect 172266 641658 172502 641894
rect 172586 641658 172822 641894
rect 172266 641338 172502 641574
rect 172586 641338 172822 641574
rect 172266 605658 172502 605894
rect 172586 605658 172822 605894
rect 172266 605338 172502 605574
rect 172586 605338 172822 605574
rect 172266 569658 172502 569894
rect 172586 569658 172822 569894
rect 172266 569338 172502 569574
rect 172586 569338 172822 569574
rect 172266 533658 172502 533894
rect 172586 533658 172822 533894
rect 172266 533338 172502 533574
rect 172586 533338 172822 533574
rect 172266 497658 172502 497894
rect 172586 497658 172822 497894
rect 172266 497338 172502 497574
rect 172586 497338 172822 497574
rect 172266 461658 172502 461894
rect 172586 461658 172822 461894
rect 172266 461338 172502 461574
rect 172586 461338 172822 461574
rect 172266 425658 172502 425894
rect 172586 425658 172822 425894
rect 172266 425338 172502 425574
rect 172586 425338 172822 425574
rect 172266 389658 172502 389894
rect 172586 389658 172822 389894
rect 172266 389338 172502 389574
rect 172586 389338 172822 389574
rect 172266 353658 172502 353894
rect 172586 353658 172822 353894
rect 172266 353338 172502 353574
rect 172586 353338 172822 353574
rect 172266 317658 172502 317894
rect 172586 317658 172822 317894
rect 172266 317338 172502 317574
rect 172586 317338 172822 317574
rect 172266 281658 172502 281894
rect 172586 281658 172822 281894
rect 172266 281338 172502 281574
rect 172586 281338 172822 281574
rect 172266 245658 172502 245894
rect 172586 245658 172822 245894
rect 172266 245338 172502 245574
rect 172586 245338 172822 245574
rect 172266 209658 172502 209894
rect 172586 209658 172822 209894
rect 172266 209338 172502 209574
rect 172586 209338 172822 209574
rect 182226 704602 182462 704838
rect 182546 704602 182782 704838
rect 182226 704282 182462 704518
rect 182546 704282 182782 704518
rect 182226 687618 182462 687854
rect 182546 687618 182782 687854
rect 182226 687298 182462 687534
rect 182546 687298 182782 687534
rect 182226 651618 182462 651854
rect 182546 651618 182782 651854
rect 182226 651298 182462 651534
rect 182546 651298 182782 651534
rect 182226 615618 182462 615854
rect 182546 615618 182782 615854
rect 182226 615298 182462 615534
rect 182546 615298 182782 615534
rect 182226 579618 182462 579854
rect 182546 579618 182782 579854
rect 182226 579298 182462 579534
rect 182546 579298 182782 579534
rect 182226 543618 182462 543854
rect 182546 543618 182782 543854
rect 182226 543298 182462 543534
rect 182546 543298 182782 543534
rect 182226 507618 182462 507854
rect 182546 507618 182782 507854
rect 182226 507298 182462 507534
rect 182546 507298 182782 507534
rect 182226 471618 182462 471854
rect 182546 471618 182782 471854
rect 182226 471298 182462 471534
rect 182546 471298 182782 471534
rect 182226 435618 182462 435854
rect 182546 435618 182782 435854
rect 182226 435298 182462 435534
rect 182546 435298 182782 435534
rect 182226 399618 182462 399854
rect 182546 399618 182782 399854
rect 182226 399298 182462 399534
rect 182546 399298 182782 399534
rect 182226 363618 182462 363854
rect 182546 363618 182782 363854
rect 182226 363298 182462 363534
rect 182546 363298 182782 363534
rect 182226 327618 182462 327854
rect 182546 327618 182782 327854
rect 182226 327298 182462 327534
rect 182546 327298 182782 327534
rect 182226 291618 182462 291854
rect 182546 291618 182782 291854
rect 182226 291298 182462 291534
rect 182546 291298 182782 291534
rect 182226 255618 182462 255854
rect 182546 255618 182782 255854
rect 182226 255298 182462 255534
rect 182546 255298 182782 255534
rect 182226 219618 182462 219854
rect 182546 219618 182782 219854
rect 182226 219298 182462 219534
rect 182546 219298 182782 219534
rect 185946 705562 186182 705798
rect 186266 705562 186502 705798
rect 185946 705242 186182 705478
rect 186266 705242 186502 705478
rect 185946 691338 186182 691574
rect 186266 691338 186502 691574
rect 185946 691018 186182 691254
rect 186266 691018 186502 691254
rect 185946 655338 186182 655574
rect 186266 655338 186502 655574
rect 185946 655018 186182 655254
rect 186266 655018 186502 655254
rect 185946 619338 186182 619574
rect 186266 619338 186502 619574
rect 185946 619018 186182 619254
rect 186266 619018 186502 619254
rect 185946 583338 186182 583574
rect 186266 583338 186502 583574
rect 185946 583018 186182 583254
rect 186266 583018 186502 583254
rect 185946 547338 186182 547574
rect 186266 547338 186502 547574
rect 185946 547018 186182 547254
rect 186266 547018 186502 547254
rect 185946 511338 186182 511574
rect 186266 511338 186502 511574
rect 185946 511018 186182 511254
rect 186266 511018 186502 511254
rect 185946 475338 186182 475574
rect 186266 475338 186502 475574
rect 185946 475018 186182 475254
rect 186266 475018 186502 475254
rect 185946 439338 186182 439574
rect 186266 439338 186502 439574
rect 185946 439018 186182 439254
rect 186266 439018 186502 439254
rect 185946 403338 186182 403574
rect 186266 403338 186502 403574
rect 185946 403018 186182 403254
rect 186266 403018 186502 403254
rect 185946 367338 186182 367574
rect 186266 367338 186502 367574
rect 185946 367018 186182 367254
rect 186266 367018 186502 367254
rect 185946 331338 186182 331574
rect 186266 331338 186502 331574
rect 185946 331018 186182 331254
rect 186266 331018 186502 331254
rect 185946 295338 186182 295574
rect 186266 295338 186502 295574
rect 185946 295018 186182 295254
rect 186266 295018 186502 295254
rect 185946 259338 186182 259574
rect 186266 259338 186502 259574
rect 185946 259018 186182 259254
rect 186266 259018 186502 259254
rect 185946 223338 186182 223574
rect 186266 223338 186502 223574
rect 185946 223018 186182 223254
rect 186266 223018 186502 223254
rect 189666 706522 189902 706758
rect 189986 706522 190222 706758
rect 189666 706202 189902 706438
rect 189986 706202 190222 706438
rect 193386 707482 193622 707718
rect 193706 707482 193942 707718
rect 193386 707162 193622 707398
rect 193706 707162 193942 707398
rect 189666 695058 189902 695294
rect 189986 695058 190222 695294
rect 189666 694738 189902 694974
rect 189986 694738 190222 694974
rect 189666 659058 189902 659294
rect 189986 659058 190222 659294
rect 189666 658738 189902 658974
rect 189986 658738 190222 658974
rect 189666 623058 189902 623294
rect 189986 623058 190222 623294
rect 189666 622738 189902 622974
rect 189986 622738 190222 622974
rect 189666 587058 189902 587294
rect 189986 587058 190222 587294
rect 189666 586738 189902 586974
rect 189986 586738 190222 586974
rect 189666 551058 189902 551294
rect 189986 551058 190222 551294
rect 189666 550738 189902 550974
rect 189986 550738 190222 550974
rect 189666 515058 189902 515294
rect 189986 515058 190222 515294
rect 189666 514738 189902 514974
rect 189986 514738 190222 514974
rect 189666 479058 189902 479294
rect 189986 479058 190222 479294
rect 189666 478738 189902 478974
rect 189986 478738 190222 478974
rect 189666 443058 189902 443294
rect 189986 443058 190222 443294
rect 189666 442738 189902 442974
rect 189986 442738 190222 442974
rect 189666 407058 189902 407294
rect 189986 407058 190222 407294
rect 189666 406738 189902 406974
rect 189986 406738 190222 406974
rect 189666 371058 189902 371294
rect 189986 371058 190222 371294
rect 189666 370738 189902 370974
rect 189986 370738 190222 370974
rect 189666 335058 189902 335294
rect 189986 335058 190222 335294
rect 189666 334738 189902 334974
rect 189986 334738 190222 334974
rect 189666 299058 189902 299294
rect 189986 299058 190222 299294
rect 189666 298738 189902 298974
rect 189986 298738 190222 298974
rect 189666 263058 189902 263294
rect 189986 263058 190222 263294
rect 189666 262738 189902 262974
rect 189986 262738 190222 262974
rect 189666 227058 189902 227294
rect 189986 227058 190222 227294
rect 189666 226738 189902 226974
rect 189986 226738 190222 226974
rect 189666 191058 189902 191294
rect 189986 191058 190222 191294
rect 189666 190738 189902 190974
rect 189986 190738 190222 190974
rect 99610 187338 99846 187574
rect 99610 187018 99846 187254
rect 130330 187338 130566 187574
rect 130330 187018 130566 187254
rect 161050 187338 161286 187574
rect 161050 187018 161286 187254
rect 114970 183618 115206 183854
rect 114970 183298 115206 183534
rect 145690 183618 145926 183854
rect 145690 183298 145926 183534
rect 176410 183618 176646 183854
rect 176410 183298 176646 183534
rect 96546 169938 96782 170174
rect 96866 169938 97102 170174
rect 96546 169618 96782 169854
rect 96866 169618 97102 169854
rect 189666 155058 189902 155294
rect 189986 155058 190222 155294
rect 189666 154738 189902 154974
rect 189986 154738 190222 154974
rect 99610 151338 99846 151574
rect 99610 151018 99846 151254
rect 130330 151338 130566 151574
rect 130330 151018 130566 151254
rect 161050 151338 161286 151574
rect 161050 151018 161286 151254
rect 114970 147618 115206 147854
rect 114970 147298 115206 147534
rect 145690 147618 145926 147854
rect 145690 147298 145926 147534
rect 176410 147618 176646 147854
rect 176410 147298 176646 147534
rect 96546 133938 96782 134174
rect 96866 133938 97102 134174
rect 96546 133618 96782 133854
rect 96866 133618 97102 133854
rect 189666 119058 189902 119294
rect 189986 119058 190222 119294
rect 189666 118738 189902 118974
rect 189986 118738 190222 118974
rect 99610 115338 99846 115574
rect 99610 115018 99846 115254
rect 130330 115338 130566 115574
rect 130330 115018 130566 115254
rect 161050 115338 161286 115574
rect 161050 115018 161286 115254
rect 114970 111618 115206 111854
rect 114970 111298 115206 111534
rect 145690 111618 145926 111854
rect 145690 111298 145926 111534
rect 176410 111618 176646 111854
rect 176410 111298 176646 111534
rect 96546 97938 96782 98174
rect 96866 97938 97102 98174
rect 96546 97618 96782 97854
rect 96866 97618 97102 97854
rect 94918 77742 95154 77978
rect 92826 58218 93062 58454
rect 93146 58218 93382 58454
rect 92826 57898 93062 58134
rect 93146 57898 93382 58134
rect 92826 22218 93062 22454
rect 93146 22218 93382 22454
rect 92826 21898 93062 22134
rect 93146 21898 93382 22134
rect 91054 4302 91290 4538
rect 89106 -4422 89342 -4186
rect 89426 -4422 89662 -4186
rect 89106 -4742 89342 -4506
rect 89426 -4742 89662 -4506
rect 96546 61938 96782 62174
rect 96866 61938 97102 62174
rect 96546 61618 96782 61854
rect 96866 61618 97102 61854
rect 96546 25938 96782 26174
rect 96866 25938 97102 26174
rect 96546 25618 96782 25854
rect 96866 25618 97102 25854
rect 92826 -5382 93062 -5146
rect 93146 -5382 93382 -5146
rect 92826 -5702 93062 -5466
rect 93146 -5702 93382 -5466
rect 100266 65658 100502 65894
rect 100586 65658 100822 65894
rect 100266 65338 100502 65574
rect 100586 65338 100822 65574
rect 100266 29658 100502 29894
rect 100586 29658 100822 29894
rect 100266 29338 100502 29574
rect 100586 29338 100822 29574
rect 96546 -6342 96782 -6106
rect 96866 -6342 97102 -6106
rect 96546 -6662 96782 -6426
rect 96866 -6662 97102 -6426
rect 100266 -7302 100502 -7066
rect 100586 -7302 100822 -7066
rect 100266 -7622 100502 -7386
rect 100586 -7622 100822 -7386
rect 110226 75618 110462 75854
rect 110546 75618 110782 75854
rect 110226 75298 110462 75534
rect 110546 75298 110782 75534
rect 110226 39618 110462 39854
rect 110546 39618 110782 39854
rect 110226 39298 110462 39534
rect 110546 39298 110782 39534
rect 113946 79338 114182 79574
rect 114266 79338 114502 79574
rect 113946 79018 114182 79254
rect 114266 79018 114502 79254
rect 113946 43338 114182 43574
rect 114266 43338 114502 43574
rect 113946 43018 114182 43254
rect 114266 43018 114502 43254
rect 113946 7338 114182 7574
rect 114266 7338 114502 7574
rect 113946 7018 114182 7254
rect 114266 7018 114502 7254
rect 117666 47058 117902 47294
rect 117986 47058 118222 47294
rect 117666 46738 117902 46974
rect 117986 46738 118222 46974
rect 117666 11058 117902 11294
rect 117986 11058 118222 11294
rect 117666 10738 117902 10974
rect 117986 10738 118222 10974
rect 113502 4302 113738 4538
rect 110226 3618 110462 3854
rect 110546 3618 110782 3854
rect 110226 3298 110462 3534
rect 110546 3298 110782 3534
rect 110226 -582 110462 -346
rect 110546 -582 110782 -346
rect 110226 -902 110462 -666
rect 110546 -902 110782 -666
rect 113946 -1542 114182 -1306
rect 114266 -1542 114502 -1306
rect 113946 -1862 114182 -1626
rect 114266 -1862 114502 -1626
rect 117666 -2502 117902 -2266
rect 117986 -2502 118222 -2266
rect 117666 -2822 117902 -2586
rect 117986 -2822 118222 -2586
rect 121386 50778 121622 51014
rect 121706 50778 121942 51014
rect 121386 50458 121622 50694
rect 121706 50458 121942 50694
rect 121386 14778 121622 15014
rect 121706 14778 121942 15014
rect 121386 14458 121622 14694
rect 121706 14458 121942 14694
rect 121386 -3462 121622 -3226
rect 121706 -3462 121942 -3226
rect 121386 -3782 121622 -3546
rect 121706 -3782 121942 -3546
rect 125106 54498 125342 54734
rect 125426 54498 125662 54734
rect 125106 54178 125342 54414
rect 125426 54178 125662 54414
rect 125106 18498 125342 18734
rect 125426 18498 125662 18734
rect 125106 18178 125342 18414
rect 125426 18178 125662 18414
rect 125106 -4422 125342 -4186
rect 125426 -4422 125662 -4186
rect 125106 -4742 125342 -4506
rect 125426 -4742 125662 -4506
rect 128826 58218 129062 58454
rect 129146 58218 129382 58454
rect 128826 57898 129062 58134
rect 129146 57898 129382 58134
rect 128826 22218 129062 22454
rect 129146 22218 129382 22454
rect 128826 21898 129062 22134
rect 129146 21898 129382 22134
rect 128826 -5382 129062 -5146
rect 129146 -5382 129382 -5146
rect 128826 -5702 129062 -5466
rect 129146 -5702 129382 -5466
rect 132546 61938 132782 62174
rect 132866 61938 133102 62174
rect 132546 61618 132782 61854
rect 132866 61618 133102 61854
rect 132546 25938 132782 26174
rect 132866 25938 133102 26174
rect 132546 25618 132782 25854
rect 132866 25618 133102 25854
rect 132546 -6342 132782 -6106
rect 132866 -6342 133102 -6106
rect 132546 -6662 132782 -6426
rect 132866 -6662 133102 -6426
rect 136266 65658 136502 65894
rect 136586 65658 136822 65894
rect 136266 65338 136502 65574
rect 136586 65338 136822 65574
rect 136266 29658 136502 29894
rect 136586 29658 136822 29894
rect 136266 29338 136502 29574
rect 136586 29338 136822 29574
rect 146226 75618 146462 75854
rect 146546 75618 146782 75854
rect 146226 75298 146462 75534
rect 146546 75298 146782 75534
rect 146226 39618 146462 39854
rect 146546 39618 146782 39854
rect 146226 39298 146462 39534
rect 146546 39298 146782 39534
rect 144966 9742 145202 9978
rect 136266 -7302 136502 -7066
rect 136586 -7302 136822 -7066
rect 136266 -7622 136502 -7386
rect 136586 -7622 136822 -7386
rect 146226 3618 146462 3854
rect 146546 3618 146782 3854
rect 146226 3298 146462 3534
rect 146546 3298 146782 3534
rect 146226 -582 146462 -346
rect 146546 -582 146782 -346
rect 146226 -902 146462 -666
rect 146546 -902 146782 -666
rect 149946 79338 150182 79574
rect 150266 79338 150502 79574
rect 149946 79018 150182 79254
rect 150266 79018 150502 79254
rect 149946 43338 150182 43574
rect 150266 43338 150502 43574
rect 149946 43018 150182 43254
rect 150266 43018 150502 43254
rect 149946 7338 150182 7574
rect 150266 7338 150502 7574
rect 149946 7018 150182 7254
rect 150266 7018 150502 7254
rect 149946 -1542 150182 -1306
rect 150266 -1542 150502 -1306
rect 149946 -1862 150182 -1626
rect 150266 -1862 150502 -1626
rect 153666 47058 153902 47294
rect 153986 47058 154222 47294
rect 153666 46738 153902 46974
rect 153986 46738 154222 46974
rect 153666 11058 153902 11294
rect 153986 11058 154222 11294
rect 153666 10738 153902 10974
rect 153986 10738 154222 10974
rect 153666 -2502 153902 -2266
rect 153986 -2502 154222 -2266
rect 153666 -2822 153902 -2586
rect 153986 -2822 154222 -2586
rect 157386 50778 157622 51014
rect 157706 50778 157942 51014
rect 157386 50458 157622 50694
rect 157706 50458 157942 50694
rect 157386 14778 157622 15014
rect 157706 14778 157942 15014
rect 157386 14458 157622 14694
rect 157706 14458 157942 14694
rect 157386 -3462 157622 -3226
rect 157706 -3462 157942 -3226
rect 157386 -3782 157622 -3546
rect 157706 -3782 157942 -3546
rect 161106 54498 161342 54734
rect 161426 54498 161662 54734
rect 161106 54178 161342 54414
rect 161426 54178 161662 54414
rect 161106 18498 161342 18734
rect 161426 18498 161662 18734
rect 161106 18178 161342 18414
rect 161426 18178 161662 18414
rect 164826 58218 165062 58454
rect 165146 58218 165382 58454
rect 164826 57898 165062 58134
rect 165146 57898 165382 58134
rect 164826 22218 165062 22454
rect 165146 22218 165382 22454
rect 164826 21898 165062 22134
rect 165146 21898 165382 22134
rect 162814 8382 163050 8618
rect 161106 -4422 161342 -4186
rect 161426 -4422 161662 -4186
rect 161106 -4742 161342 -4506
rect 161426 -4742 161662 -4506
rect 164826 -5382 165062 -5146
rect 165146 -5382 165382 -5146
rect 164826 -5702 165062 -5466
rect 165146 -5702 165382 -5466
rect 168546 61938 168782 62174
rect 168866 61938 169102 62174
rect 168546 61618 168782 61854
rect 168866 61618 169102 61854
rect 168546 25938 168782 26174
rect 168866 25938 169102 26174
rect 168546 25618 168782 25854
rect 168866 25618 169102 25854
rect 168546 -6342 168782 -6106
rect 168866 -6342 169102 -6106
rect 168546 -6662 168782 -6426
rect 168866 -6662 169102 -6426
rect 175142 77892 175378 77978
rect 175142 77828 175228 77892
rect 175228 77828 175292 77892
rect 175292 77828 175378 77892
rect 175142 77742 175378 77828
rect 177166 77742 177402 77978
rect 172266 65658 172502 65894
rect 172586 65658 172822 65894
rect 172266 65338 172502 65574
rect 172586 65338 172822 65574
rect 172266 29658 172502 29894
rect 172586 29658 172822 29894
rect 172266 29338 172502 29574
rect 172586 29338 172822 29574
rect 182226 75618 182462 75854
rect 182546 75618 182782 75854
rect 182226 75298 182462 75534
rect 182546 75298 182782 75534
rect 182226 39618 182462 39854
rect 182546 39618 182782 39854
rect 182226 39298 182462 39534
rect 182546 39298 182782 39534
rect 172266 -7302 172502 -7066
rect 172586 -7302 172822 -7066
rect 172266 -7622 172502 -7386
rect 172586 -7622 172822 -7386
rect 182226 3618 182462 3854
rect 182546 3618 182782 3854
rect 182226 3298 182462 3534
rect 182546 3298 182782 3534
rect 182226 -582 182462 -346
rect 182546 -582 182782 -346
rect 182226 -902 182462 -666
rect 182546 -902 182782 -666
rect 185946 79338 186182 79574
rect 186266 79338 186502 79574
rect 185946 79018 186182 79254
rect 186266 79018 186502 79254
rect 185946 43338 186182 43574
rect 186266 43338 186502 43574
rect 185946 43018 186182 43254
rect 186266 43018 186502 43254
rect 185946 7338 186182 7574
rect 186266 7338 186502 7574
rect 185946 7018 186182 7254
rect 186266 7018 186502 7254
rect 189666 83058 189902 83294
rect 189986 83058 190222 83294
rect 189666 82738 189902 82974
rect 189986 82738 190222 82974
rect 189666 47058 189902 47294
rect 189986 47058 190222 47294
rect 189666 46738 189902 46974
rect 189986 46738 190222 46974
rect 189666 11058 189902 11294
rect 189986 11058 190222 11294
rect 189666 10738 189902 10974
rect 189986 10738 190222 10974
rect 185946 -1542 186182 -1306
rect 186266 -1542 186502 -1306
rect 185946 -1862 186182 -1626
rect 186266 -1862 186502 -1626
rect 190598 5662 190834 5898
rect 191334 11782 191570 12018
rect 193386 698778 193622 699014
rect 193706 698778 193942 699014
rect 193386 698458 193622 698694
rect 193706 698458 193942 698694
rect 193386 662778 193622 663014
rect 193706 662778 193942 663014
rect 193386 662458 193622 662694
rect 193706 662458 193942 662694
rect 193386 626778 193622 627014
rect 193706 626778 193942 627014
rect 193386 626458 193622 626694
rect 193706 626458 193942 626694
rect 193386 590778 193622 591014
rect 193706 590778 193942 591014
rect 193386 590458 193622 590694
rect 193706 590458 193942 590694
rect 193386 554778 193622 555014
rect 193706 554778 193942 555014
rect 193386 554458 193622 554694
rect 193706 554458 193942 554694
rect 193386 518778 193622 519014
rect 193706 518778 193942 519014
rect 193386 518458 193622 518694
rect 193706 518458 193942 518694
rect 193386 482778 193622 483014
rect 193706 482778 193942 483014
rect 193386 482458 193622 482694
rect 193706 482458 193942 482694
rect 193386 446778 193622 447014
rect 193706 446778 193942 447014
rect 193386 446458 193622 446694
rect 193706 446458 193942 446694
rect 193386 410778 193622 411014
rect 193706 410778 193942 411014
rect 193386 410458 193622 410694
rect 193706 410458 193942 410694
rect 193386 374778 193622 375014
rect 193706 374778 193942 375014
rect 193386 374458 193622 374694
rect 193706 374458 193942 374694
rect 193386 338778 193622 339014
rect 193706 338778 193942 339014
rect 193386 338458 193622 338694
rect 193706 338458 193942 338694
rect 193386 302778 193622 303014
rect 193706 302778 193942 303014
rect 193386 302458 193622 302694
rect 193706 302458 193942 302694
rect 193386 266778 193622 267014
rect 193706 266778 193942 267014
rect 193386 266458 193622 266694
rect 193706 266458 193942 266694
rect 193386 230778 193622 231014
rect 193706 230778 193942 231014
rect 193386 230458 193622 230694
rect 193706 230458 193942 230694
rect 193386 194778 193622 195014
rect 193706 194778 193942 195014
rect 193386 194458 193622 194694
rect 193706 194458 193942 194694
rect 193386 158778 193622 159014
rect 193706 158778 193942 159014
rect 193386 158458 193622 158694
rect 193706 158458 193942 158694
rect 193386 122778 193622 123014
rect 193706 122778 193942 123014
rect 193386 122458 193622 122694
rect 193706 122458 193942 122694
rect 193386 86778 193622 87014
rect 193706 86778 193942 87014
rect 193386 86458 193622 86694
rect 193706 86458 193942 86694
rect 193386 50778 193622 51014
rect 193706 50778 193942 51014
rect 193386 50458 193622 50694
rect 193706 50458 193942 50694
rect 191702 6342 191938 6578
rect 193386 14778 193622 15014
rect 193706 14778 193942 15014
rect 193386 14458 193622 14694
rect 193706 14458 193942 14694
rect 191334 4982 191570 5218
rect 189666 -2502 189902 -2266
rect 189986 -2502 190222 -2266
rect 189666 -2822 189902 -2586
rect 189986 -2822 190222 -2586
rect 193386 -3462 193622 -3226
rect 193706 -3462 193942 -3226
rect 193386 -3782 193622 -3546
rect 193706 -3782 193942 -3546
rect 197106 708442 197342 708678
rect 197426 708442 197662 708678
rect 197106 708122 197342 708358
rect 197426 708122 197662 708358
rect 197106 666498 197342 666734
rect 197426 666498 197662 666734
rect 197106 666178 197342 666414
rect 197426 666178 197662 666414
rect 197106 630498 197342 630734
rect 197426 630498 197662 630734
rect 197106 630178 197342 630414
rect 197426 630178 197662 630414
rect 197106 594498 197342 594734
rect 197426 594498 197662 594734
rect 197106 594178 197342 594414
rect 197426 594178 197662 594414
rect 197106 558498 197342 558734
rect 197426 558498 197662 558734
rect 197106 558178 197342 558414
rect 197426 558178 197662 558414
rect 197106 522498 197342 522734
rect 197426 522498 197662 522734
rect 197106 522178 197342 522414
rect 197426 522178 197662 522414
rect 197106 486498 197342 486734
rect 197426 486498 197662 486734
rect 197106 486178 197342 486414
rect 197426 486178 197662 486414
rect 197106 450498 197342 450734
rect 197426 450498 197662 450734
rect 197106 450178 197342 450414
rect 197426 450178 197662 450414
rect 197106 414498 197342 414734
rect 197426 414498 197662 414734
rect 197106 414178 197342 414414
rect 197426 414178 197662 414414
rect 197106 378498 197342 378734
rect 197426 378498 197662 378734
rect 197106 378178 197342 378414
rect 197426 378178 197662 378414
rect 197106 342498 197342 342734
rect 197426 342498 197662 342734
rect 197106 342178 197342 342414
rect 197426 342178 197662 342414
rect 197106 306498 197342 306734
rect 197426 306498 197662 306734
rect 197106 306178 197342 306414
rect 197426 306178 197662 306414
rect 197106 270498 197342 270734
rect 197426 270498 197662 270734
rect 197106 270178 197342 270414
rect 197426 270178 197662 270414
rect 197106 234498 197342 234734
rect 197426 234498 197662 234734
rect 197106 234178 197342 234414
rect 197426 234178 197662 234414
rect 197106 198498 197342 198734
rect 197426 198498 197662 198734
rect 197106 198178 197342 198414
rect 197426 198178 197662 198414
rect 197106 162498 197342 162734
rect 197426 162498 197662 162734
rect 197106 162178 197342 162414
rect 197426 162178 197662 162414
rect 197106 126498 197342 126734
rect 197426 126498 197662 126734
rect 197106 126178 197342 126414
rect 197426 126178 197662 126414
rect 197106 90498 197342 90734
rect 197426 90498 197662 90734
rect 197106 90178 197342 90414
rect 197426 90178 197662 90414
rect 197106 54498 197342 54734
rect 197426 54498 197662 54734
rect 197106 54178 197342 54414
rect 197426 54178 197662 54414
rect 197106 18498 197342 18734
rect 197426 18498 197662 18734
rect 197106 18178 197342 18414
rect 197426 18178 197662 18414
rect 197106 -4422 197342 -4186
rect 197426 -4422 197662 -4186
rect 197106 -4742 197342 -4506
rect 197426 -4742 197662 -4506
rect 200826 709402 201062 709638
rect 201146 709402 201382 709638
rect 200826 709082 201062 709318
rect 201146 709082 201382 709318
rect 200826 670218 201062 670454
rect 201146 670218 201382 670454
rect 200826 669898 201062 670134
rect 201146 669898 201382 670134
rect 200826 634218 201062 634454
rect 201146 634218 201382 634454
rect 200826 633898 201062 634134
rect 201146 633898 201382 634134
rect 200826 598218 201062 598454
rect 201146 598218 201382 598454
rect 200826 597898 201062 598134
rect 201146 597898 201382 598134
rect 200826 562218 201062 562454
rect 201146 562218 201382 562454
rect 200826 561898 201062 562134
rect 201146 561898 201382 562134
rect 200826 526218 201062 526454
rect 201146 526218 201382 526454
rect 200826 525898 201062 526134
rect 201146 525898 201382 526134
rect 200826 490218 201062 490454
rect 201146 490218 201382 490454
rect 200826 489898 201062 490134
rect 201146 489898 201382 490134
rect 200826 454218 201062 454454
rect 201146 454218 201382 454454
rect 200826 453898 201062 454134
rect 201146 453898 201382 454134
rect 200826 418218 201062 418454
rect 201146 418218 201382 418454
rect 200826 417898 201062 418134
rect 201146 417898 201382 418134
rect 200826 382218 201062 382454
rect 201146 382218 201382 382454
rect 200826 381898 201062 382134
rect 201146 381898 201382 382134
rect 200826 346218 201062 346454
rect 201146 346218 201382 346454
rect 200826 345898 201062 346134
rect 201146 345898 201382 346134
rect 200826 310218 201062 310454
rect 201146 310218 201382 310454
rect 200826 309898 201062 310134
rect 201146 309898 201382 310134
rect 200826 274218 201062 274454
rect 201146 274218 201382 274454
rect 200826 273898 201062 274134
rect 201146 273898 201382 274134
rect 200826 238218 201062 238454
rect 201146 238218 201382 238454
rect 200826 237898 201062 238134
rect 201146 237898 201382 238134
rect 200826 202218 201062 202454
rect 201146 202218 201382 202454
rect 200826 201898 201062 202134
rect 201146 201898 201382 202134
rect 200826 166218 201062 166454
rect 201146 166218 201382 166454
rect 200826 165898 201062 166134
rect 201146 165898 201382 166134
rect 200826 130218 201062 130454
rect 201146 130218 201382 130454
rect 200826 129898 201062 130134
rect 201146 129898 201382 130134
rect 200826 94218 201062 94454
rect 201146 94218 201382 94454
rect 200826 93898 201062 94134
rect 201146 93898 201382 94134
rect 200826 58218 201062 58454
rect 201146 58218 201382 58454
rect 200826 57898 201062 58134
rect 201146 57898 201382 58134
rect 200826 22218 201062 22454
rect 201146 22218 201382 22454
rect 200826 21898 201062 22134
rect 201146 21898 201382 22134
rect 204546 710362 204782 710598
rect 204866 710362 205102 710598
rect 204546 710042 204782 710278
rect 204866 710042 205102 710278
rect 204546 673938 204782 674174
rect 204866 673938 205102 674174
rect 204546 673618 204782 673854
rect 204866 673618 205102 673854
rect 204546 637938 204782 638174
rect 204866 637938 205102 638174
rect 204546 637618 204782 637854
rect 204866 637618 205102 637854
rect 204546 601938 204782 602174
rect 204866 601938 205102 602174
rect 204546 601618 204782 601854
rect 204866 601618 205102 601854
rect 204546 565938 204782 566174
rect 204866 565938 205102 566174
rect 204546 565618 204782 565854
rect 204866 565618 205102 565854
rect 204546 529938 204782 530174
rect 204866 529938 205102 530174
rect 204546 529618 204782 529854
rect 204866 529618 205102 529854
rect 204546 493938 204782 494174
rect 204866 493938 205102 494174
rect 204546 493618 204782 493854
rect 204866 493618 205102 493854
rect 204546 457938 204782 458174
rect 204866 457938 205102 458174
rect 204546 457618 204782 457854
rect 204866 457618 205102 457854
rect 204546 421938 204782 422174
rect 204866 421938 205102 422174
rect 204546 421618 204782 421854
rect 204866 421618 205102 421854
rect 204546 385938 204782 386174
rect 204866 385938 205102 386174
rect 204546 385618 204782 385854
rect 204866 385618 205102 385854
rect 204546 349938 204782 350174
rect 204866 349938 205102 350174
rect 204546 349618 204782 349854
rect 204866 349618 205102 349854
rect 204546 313938 204782 314174
rect 204866 313938 205102 314174
rect 204546 313618 204782 313854
rect 204866 313618 205102 313854
rect 204546 277938 204782 278174
rect 204866 277938 205102 278174
rect 204546 277618 204782 277854
rect 204866 277618 205102 277854
rect 204546 241938 204782 242174
rect 204866 241938 205102 242174
rect 204546 241618 204782 241854
rect 204866 241618 205102 241854
rect 204546 205938 204782 206174
rect 204866 205938 205102 206174
rect 204546 205618 204782 205854
rect 204866 205618 205102 205854
rect 204546 169938 204782 170174
rect 204866 169938 205102 170174
rect 204546 169618 204782 169854
rect 204866 169618 205102 169854
rect 204546 133938 204782 134174
rect 204866 133938 205102 134174
rect 204546 133618 204782 133854
rect 204866 133618 205102 133854
rect 204546 97938 204782 98174
rect 204866 97938 205102 98174
rect 204546 97618 204782 97854
rect 204866 97618 205102 97854
rect 204546 61938 204782 62174
rect 204866 61938 205102 62174
rect 204546 61618 204782 61854
rect 204866 61618 205102 61854
rect 204546 25938 204782 26174
rect 204866 25938 205102 26174
rect 204546 25618 204782 25854
rect 204866 25618 205102 25854
rect 204030 4302 204266 4538
rect 200826 -5382 201062 -5146
rect 201146 -5382 201382 -5146
rect 200826 -5702 201062 -5466
rect 201146 -5702 201382 -5466
rect 204546 -6342 204782 -6106
rect 204866 -6342 205102 -6106
rect 204546 -6662 204782 -6426
rect 204866 -6662 205102 -6426
rect 208266 711322 208502 711558
rect 208586 711322 208822 711558
rect 208266 711002 208502 711238
rect 208586 711002 208822 711238
rect 208266 677658 208502 677894
rect 208586 677658 208822 677894
rect 208266 677338 208502 677574
rect 208586 677338 208822 677574
rect 208266 641658 208502 641894
rect 208586 641658 208822 641894
rect 208266 641338 208502 641574
rect 208586 641338 208822 641574
rect 208266 605658 208502 605894
rect 208586 605658 208822 605894
rect 208266 605338 208502 605574
rect 208586 605338 208822 605574
rect 208266 569658 208502 569894
rect 208586 569658 208822 569894
rect 208266 569338 208502 569574
rect 208586 569338 208822 569574
rect 208266 533658 208502 533894
rect 208586 533658 208822 533894
rect 208266 533338 208502 533574
rect 208586 533338 208822 533574
rect 208266 497658 208502 497894
rect 208586 497658 208822 497894
rect 208266 497338 208502 497574
rect 208586 497338 208822 497574
rect 208266 461658 208502 461894
rect 208586 461658 208822 461894
rect 208266 461338 208502 461574
rect 208586 461338 208822 461574
rect 208266 425658 208502 425894
rect 208586 425658 208822 425894
rect 208266 425338 208502 425574
rect 208586 425338 208822 425574
rect 208266 389658 208502 389894
rect 208586 389658 208822 389894
rect 208266 389338 208502 389574
rect 208586 389338 208822 389574
rect 208266 353658 208502 353894
rect 208586 353658 208822 353894
rect 208266 353338 208502 353574
rect 208586 353338 208822 353574
rect 208266 317658 208502 317894
rect 208586 317658 208822 317894
rect 208266 317338 208502 317574
rect 208586 317338 208822 317574
rect 208266 281658 208502 281894
rect 208586 281658 208822 281894
rect 208266 281338 208502 281574
rect 208586 281338 208822 281574
rect 208266 245658 208502 245894
rect 208586 245658 208822 245894
rect 208266 245338 208502 245574
rect 208586 245338 208822 245574
rect 208266 209658 208502 209894
rect 208586 209658 208822 209894
rect 208266 209338 208502 209574
rect 208586 209338 208822 209574
rect 208266 173658 208502 173894
rect 208586 173658 208822 173894
rect 208266 173338 208502 173574
rect 208586 173338 208822 173574
rect 208266 137658 208502 137894
rect 208586 137658 208822 137894
rect 208266 137338 208502 137574
rect 208586 137338 208822 137574
rect 208266 101658 208502 101894
rect 208586 101658 208822 101894
rect 208266 101338 208502 101574
rect 208586 101338 208822 101574
rect 208266 65658 208502 65894
rect 208586 65658 208822 65894
rect 208266 65338 208502 65574
rect 208586 65338 208822 65574
rect 208266 29658 208502 29894
rect 208586 29658 208822 29894
rect 208266 29338 208502 29574
rect 208586 29338 208822 29574
rect 218226 704602 218462 704838
rect 218546 704602 218782 704838
rect 218226 704282 218462 704518
rect 218546 704282 218782 704518
rect 218226 687618 218462 687854
rect 218546 687618 218782 687854
rect 218226 687298 218462 687534
rect 218546 687298 218782 687534
rect 218226 651618 218462 651854
rect 218546 651618 218782 651854
rect 218226 651298 218462 651534
rect 218546 651298 218782 651534
rect 218226 615618 218462 615854
rect 218546 615618 218782 615854
rect 218226 615298 218462 615534
rect 218546 615298 218782 615534
rect 218226 579618 218462 579854
rect 218546 579618 218782 579854
rect 218226 579298 218462 579534
rect 218546 579298 218782 579534
rect 218226 543618 218462 543854
rect 218546 543618 218782 543854
rect 218226 543298 218462 543534
rect 218546 543298 218782 543534
rect 218226 507618 218462 507854
rect 218546 507618 218782 507854
rect 218226 507298 218462 507534
rect 218546 507298 218782 507534
rect 218226 471618 218462 471854
rect 218546 471618 218782 471854
rect 218226 471298 218462 471534
rect 218546 471298 218782 471534
rect 218226 435618 218462 435854
rect 218546 435618 218782 435854
rect 218226 435298 218462 435534
rect 218546 435298 218782 435534
rect 218226 399618 218462 399854
rect 218546 399618 218782 399854
rect 218226 399298 218462 399534
rect 218546 399298 218782 399534
rect 218226 363618 218462 363854
rect 218546 363618 218782 363854
rect 218226 363298 218462 363534
rect 218546 363298 218782 363534
rect 218226 327618 218462 327854
rect 218546 327618 218782 327854
rect 218226 327298 218462 327534
rect 218546 327298 218782 327534
rect 218226 291618 218462 291854
rect 218546 291618 218782 291854
rect 218226 291298 218462 291534
rect 218546 291298 218782 291534
rect 218226 255618 218462 255854
rect 218546 255618 218782 255854
rect 218226 255298 218462 255534
rect 218546 255298 218782 255534
rect 218226 219618 218462 219854
rect 218546 219618 218782 219854
rect 218226 219298 218462 219534
rect 218546 219298 218782 219534
rect 218226 183618 218462 183854
rect 218546 183618 218782 183854
rect 218226 183298 218462 183534
rect 218546 183298 218782 183534
rect 218226 147618 218462 147854
rect 218546 147618 218782 147854
rect 218226 147298 218462 147534
rect 218546 147298 218782 147534
rect 218226 111618 218462 111854
rect 218546 111618 218782 111854
rect 218226 111298 218462 111534
rect 218546 111298 218782 111534
rect 218226 75618 218462 75854
rect 218546 75618 218782 75854
rect 218226 75298 218462 75534
rect 218546 75298 218782 75534
rect 218226 39618 218462 39854
rect 218546 39618 218782 39854
rect 218226 39298 218462 39534
rect 218546 39298 218782 39534
rect 208266 -7302 208502 -7066
rect 208586 -7302 208822 -7066
rect 208266 -7622 208502 -7386
rect 208586 -7622 208822 -7386
rect 218226 3618 218462 3854
rect 218546 3618 218782 3854
rect 218226 3298 218462 3534
rect 218546 3298 218782 3534
rect 218226 -582 218462 -346
rect 218546 -582 218782 -346
rect 218226 -902 218462 -666
rect 218546 -902 218782 -666
rect 221946 705562 222182 705798
rect 222266 705562 222502 705798
rect 221946 705242 222182 705478
rect 222266 705242 222502 705478
rect 221946 691338 222182 691574
rect 222266 691338 222502 691574
rect 221946 691018 222182 691254
rect 222266 691018 222502 691254
rect 221946 655338 222182 655574
rect 222266 655338 222502 655574
rect 221946 655018 222182 655254
rect 222266 655018 222502 655254
rect 221946 619338 222182 619574
rect 222266 619338 222502 619574
rect 221946 619018 222182 619254
rect 222266 619018 222502 619254
rect 221946 583338 222182 583574
rect 222266 583338 222502 583574
rect 221946 583018 222182 583254
rect 222266 583018 222502 583254
rect 221946 547338 222182 547574
rect 222266 547338 222502 547574
rect 221946 547018 222182 547254
rect 222266 547018 222502 547254
rect 221946 511338 222182 511574
rect 222266 511338 222502 511574
rect 221946 511018 222182 511254
rect 222266 511018 222502 511254
rect 221946 475338 222182 475574
rect 222266 475338 222502 475574
rect 221946 475018 222182 475254
rect 222266 475018 222502 475254
rect 221946 439338 222182 439574
rect 222266 439338 222502 439574
rect 221946 439018 222182 439254
rect 222266 439018 222502 439254
rect 221946 403338 222182 403574
rect 222266 403338 222502 403574
rect 221946 403018 222182 403254
rect 222266 403018 222502 403254
rect 221946 367338 222182 367574
rect 222266 367338 222502 367574
rect 221946 367018 222182 367254
rect 222266 367018 222502 367254
rect 221946 331338 222182 331574
rect 222266 331338 222502 331574
rect 221946 331018 222182 331254
rect 222266 331018 222502 331254
rect 221946 295338 222182 295574
rect 222266 295338 222502 295574
rect 221946 295018 222182 295254
rect 222266 295018 222502 295254
rect 221946 259338 222182 259574
rect 222266 259338 222502 259574
rect 221946 259018 222182 259254
rect 222266 259018 222502 259254
rect 221946 223338 222182 223574
rect 222266 223338 222502 223574
rect 221946 223018 222182 223254
rect 222266 223018 222502 223254
rect 221946 187338 222182 187574
rect 222266 187338 222502 187574
rect 221946 187018 222182 187254
rect 222266 187018 222502 187254
rect 221946 151338 222182 151574
rect 222266 151338 222502 151574
rect 221946 151018 222182 151254
rect 222266 151018 222502 151254
rect 221946 115338 222182 115574
rect 222266 115338 222502 115574
rect 221946 115018 222182 115254
rect 222266 115018 222502 115254
rect 221946 79338 222182 79574
rect 222266 79338 222502 79574
rect 221946 79018 222182 79254
rect 222266 79018 222502 79254
rect 221946 43338 222182 43574
rect 222266 43338 222502 43574
rect 221946 43018 222182 43254
rect 222266 43018 222502 43254
rect 221946 7338 222182 7574
rect 222266 7338 222502 7574
rect 221946 7018 222182 7254
rect 222266 7018 222502 7254
rect 221946 -1542 222182 -1306
rect 222266 -1542 222502 -1306
rect 221946 -1862 222182 -1626
rect 222266 -1862 222502 -1626
rect 225666 706522 225902 706758
rect 225986 706522 226222 706758
rect 225666 706202 225902 706438
rect 225986 706202 226222 706438
rect 225666 695058 225902 695294
rect 225986 695058 226222 695294
rect 225666 694738 225902 694974
rect 225986 694738 226222 694974
rect 225666 659058 225902 659294
rect 225986 659058 226222 659294
rect 225666 658738 225902 658974
rect 225986 658738 226222 658974
rect 225666 623058 225902 623294
rect 225986 623058 226222 623294
rect 225666 622738 225902 622974
rect 225986 622738 226222 622974
rect 225666 587058 225902 587294
rect 225986 587058 226222 587294
rect 225666 586738 225902 586974
rect 225986 586738 226222 586974
rect 225666 551058 225902 551294
rect 225986 551058 226222 551294
rect 225666 550738 225902 550974
rect 225986 550738 226222 550974
rect 225666 515058 225902 515294
rect 225986 515058 226222 515294
rect 225666 514738 225902 514974
rect 225986 514738 226222 514974
rect 225666 479058 225902 479294
rect 225986 479058 226222 479294
rect 225666 478738 225902 478974
rect 225986 478738 226222 478974
rect 225666 443058 225902 443294
rect 225986 443058 226222 443294
rect 225666 442738 225902 442974
rect 225986 442738 226222 442974
rect 225666 407058 225902 407294
rect 225986 407058 226222 407294
rect 225666 406738 225902 406974
rect 225986 406738 226222 406974
rect 225666 371058 225902 371294
rect 225986 371058 226222 371294
rect 225666 370738 225902 370974
rect 225986 370738 226222 370974
rect 225666 335058 225902 335294
rect 225986 335058 226222 335294
rect 225666 334738 225902 334974
rect 225986 334738 226222 334974
rect 225666 299058 225902 299294
rect 225986 299058 226222 299294
rect 225666 298738 225902 298974
rect 225986 298738 226222 298974
rect 225666 263058 225902 263294
rect 225986 263058 226222 263294
rect 225666 262738 225902 262974
rect 225986 262738 226222 262974
rect 225666 227058 225902 227294
rect 225986 227058 226222 227294
rect 225666 226738 225902 226974
rect 225986 226738 226222 226974
rect 225666 191058 225902 191294
rect 225986 191058 226222 191294
rect 225666 190738 225902 190974
rect 225986 190738 226222 190974
rect 225666 155058 225902 155294
rect 225986 155058 226222 155294
rect 225666 154738 225902 154974
rect 225986 154738 226222 154974
rect 225666 119058 225902 119294
rect 225986 119058 226222 119294
rect 225666 118738 225902 118974
rect 225986 118738 226222 118974
rect 225666 83058 225902 83294
rect 225986 83058 226222 83294
rect 225666 82738 225902 82974
rect 225986 82738 226222 82974
rect 225666 47058 225902 47294
rect 225986 47058 226222 47294
rect 225666 46738 225902 46974
rect 225986 46738 226222 46974
rect 225666 11058 225902 11294
rect 225986 11058 226222 11294
rect 225666 10738 225902 10974
rect 225986 10738 226222 10974
rect 225666 -2502 225902 -2266
rect 225986 -2502 226222 -2266
rect 225666 -2822 225902 -2586
rect 225986 -2822 226222 -2586
rect 229386 707482 229622 707718
rect 229706 707482 229942 707718
rect 229386 707162 229622 707398
rect 229706 707162 229942 707398
rect 229386 698778 229622 699014
rect 229706 698778 229942 699014
rect 229386 698458 229622 698694
rect 229706 698458 229942 698694
rect 229386 662778 229622 663014
rect 229706 662778 229942 663014
rect 229386 662458 229622 662694
rect 229706 662458 229942 662694
rect 229386 626778 229622 627014
rect 229706 626778 229942 627014
rect 229386 626458 229622 626694
rect 229706 626458 229942 626694
rect 229386 590778 229622 591014
rect 229706 590778 229942 591014
rect 229386 590458 229622 590694
rect 229706 590458 229942 590694
rect 229386 554778 229622 555014
rect 229706 554778 229942 555014
rect 229386 554458 229622 554694
rect 229706 554458 229942 554694
rect 229386 518778 229622 519014
rect 229706 518778 229942 519014
rect 229386 518458 229622 518694
rect 229706 518458 229942 518694
rect 229386 482778 229622 483014
rect 229706 482778 229942 483014
rect 229386 482458 229622 482694
rect 229706 482458 229942 482694
rect 229386 446778 229622 447014
rect 229706 446778 229942 447014
rect 229386 446458 229622 446694
rect 229706 446458 229942 446694
rect 229386 410778 229622 411014
rect 229706 410778 229942 411014
rect 229386 410458 229622 410694
rect 229706 410458 229942 410694
rect 229386 374778 229622 375014
rect 229706 374778 229942 375014
rect 229386 374458 229622 374694
rect 229706 374458 229942 374694
rect 229386 338778 229622 339014
rect 229706 338778 229942 339014
rect 229386 338458 229622 338694
rect 229706 338458 229942 338694
rect 229386 302778 229622 303014
rect 229706 302778 229942 303014
rect 229386 302458 229622 302694
rect 229706 302458 229942 302694
rect 229386 266778 229622 267014
rect 229706 266778 229942 267014
rect 229386 266458 229622 266694
rect 229706 266458 229942 266694
rect 229386 230778 229622 231014
rect 229706 230778 229942 231014
rect 229386 230458 229622 230694
rect 229706 230458 229942 230694
rect 229386 194778 229622 195014
rect 229706 194778 229942 195014
rect 229386 194458 229622 194694
rect 229706 194458 229942 194694
rect 229386 158778 229622 159014
rect 229706 158778 229942 159014
rect 229386 158458 229622 158694
rect 229706 158458 229942 158694
rect 229386 122778 229622 123014
rect 229706 122778 229942 123014
rect 229386 122458 229622 122694
rect 229706 122458 229942 122694
rect 229386 86778 229622 87014
rect 229706 86778 229942 87014
rect 229386 86458 229622 86694
rect 229706 86458 229942 86694
rect 229386 50778 229622 51014
rect 229706 50778 229942 51014
rect 229386 50458 229622 50694
rect 229706 50458 229942 50694
rect 229386 14778 229622 15014
rect 229706 14778 229942 15014
rect 229386 14458 229622 14694
rect 229706 14458 229942 14694
rect 229386 -3462 229622 -3226
rect 229706 -3462 229942 -3226
rect 229386 -3782 229622 -3546
rect 229706 -3782 229942 -3546
rect 233106 708442 233342 708678
rect 233426 708442 233662 708678
rect 233106 708122 233342 708358
rect 233426 708122 233662 708358
rect 233106 666498 233342 666734
rect 233426 666498 233662 666734
rect 233106 666178 233342 666414
rect 233426 666178 233662 666414
rect 233106 630498 233342 630734
rect 233426 630498 233662 630734
rect 233106 630178 233342 630414
rect 233426 630178 233662 630414
rect 233106 594498 233342 594734
rect 233426 594498 233662 594734
rect 233106 594178 233342 594414
rect 233426 594178 233662 594414
rect 233106 558498 233342 558734
rect 233426 558498 233662 558734
rect 233106 558178 233342 558414
rect 233426 558178 233662 558414
rect 233106 522498 233342 522734
rect 233426 522498 233662 522734
rect 233106 522178 233342 522414
rect 233426 522178 233662 522414
rect 233106 486498 233342 486734
rect 233426 486498 233662 486734
rect 233106 486178 233342 486414
rect 233426 486178 233662 486414
rect 233106 450498 233342 450734
rect 233426 450498 233662 450734
rect 233106 450178 233342 450414
rect 233426 450178 233662 450414
rect 233106 414498 233342 414734
rect 233426 414498 233662 414734
rect 233106 414178 233342 414414
rect 233426 414178 233662 414414
rect 233106 378498 233342 378734
rect 233426 378498 233662 378734
rect 233106 378178 233342 378414
rect 233426 378178 233662 378414
rect 233106 342498 233342 342734
rect 233426 342498 233662 342734
rect 233106 342178 233342 342414
rect 233426 342178 233662 342414
rect 233106 306498 233342 306734
rect 233426 306498 233662 306734
rect 233106 306178 233342 306414
rect 233426 306178 233662 306414
rect 233106 270498 233342 270734
rect 233426 270498 233662 270734
rect 233106 270178 233342 270414
rect 233426 270178 233662 270414
rect 233106 234498 233342 234734
rect 233426 234498 233662 234734
rect 233106 234178 233342 234414
rect 233426 234178 233662 234414
rect 233106 198498 233342 198734
rect 233426 198498 233662 198734
rect 233106 198178 233342 198414
rect 233426 198178 233662 198414
rect 233106 162498 233342 162734
rect 233426 162498 233662 162734
rect 233106 162178 233342 162414
rect 233426 162178 233662 162414
rect 233106 126498 233342 126734
rect 233426 126498 233662 126734
rect 233106 126178 233342 126414
rect 233426 126178 233662 126414
rect 233106 90498 233342 90734
rect 233426 90498 233662 90734
rect 233106 90178 233342 90414
rect 233426 90178 233662 90414
rect 233106 54498 233342 54734
rect 233426 54498 233662 54734
rect 233106 54178 233342 54414
rect 233426 54178 233662 54414
rect 233106 18498 233342 18734
rect 233426 18498 233662 18734
rect 233106 18178 233342 18414
rect 233426 18178 233662 18414
rect 233106 -4422 233342 -4186
rect 233426 -4422 233662 -4186
rect 233106 -4742 233342 -4506
rect 233426 -4742 233662 -4506
rect 236826 709402 237062 709638
rect 237146 709402 237382 709638
rect 236826 709082 237062 709318
rect 237146 709082 237382 709318
rect 236826 670218 237062 670454
rect 237146 670218 237382 670454
rect 236826 669898 237062 670134
rect 237146 669898 237382 670134
rect 236826 634218 237062 634454
rect 237146 634218 237382 634454
rect 236826 633898 237062 634134
rect 237146 633898 237382 634134
rect 236826 598218 237062 598454
rect 237146 598218 237382 598454
rect 236826 597898 237062 598134
rect 237146 597898 237382 598134
rect 236826 562218 237062 562454
rect 237146 562218 237382 562454
rect 236826 561898 237062 562134
rect 237146 561898 237382 562134
rect 236826 526218 237062 526454
rect 237146 526218 237382 526454
rect 236826 525898 237062 526134
rect 237146 525898 237382 526134
rect 236826 490218 237062 490454
rect 237146 490218 237382 490454
rect 236826 489898 237062 490134
rect 237146 489898 237382 490134
rect 236826 454218 237062 454454
rect 237146 454218 237382 454454
rect 236826 453898 237062 454134
rect 237146 453898 237382 454134
rect 236826 418218 237062 418454
rect 237146 418218 237382 418454
rect 236826 417898 237062 418134
rect 237146 417898 237382 418134
rect 236826 382218 237062 382454
rect 237146 382218 237382 382454
rect 236826 381898 237062 382134
rect 237146 381898 237382 382134
rect 236826 346218 237062 346454
rect 237146 346218 237382 346454
rect 236826 345898 237062 346134
rect 237146 345898 237382 346134
rect 236826 310218 237062 310454
rect 237146 310218 237382 310454
rect 236826 309898 237062 310134
rect 237146 309898 237382 310134
rect 236826 274218 237062 274454
rect 237146 274218 237382 274454
rect 236826 273898 237062 274134
rect 237146 273898 237382 274134
rect 236826 238218 237062 238454
rect 237146 238218 237382 238454
rect 236826 237898 237062 238134
rect 237146 237898 237382 238134
rect 236826 202218 237062 202454
rect 237146 202218 237382 202454
rect 236826 201898 237062 202134
rect 237146 201898 237382 202134
rect 236826 166218 237062 166454
rect 237146 166218 237382 166454
rect 236826 165898 237062 166134
rect 237146 165898 237382 166134
rect 236826 130218 237062 130454
rect 237146 130218 237382 130454
rect 236826 129898 237062 130134
rect 237146 129898 237382 130134
rect 236826 94218 237062 94454
rect 237146 94218 237382 94454
rect 236826 93898 237062 94134
rect 237146 93898 237382 94134
rect 236826 58218 237062 58454
rect 237146 58218 237382 58454
rect 236826 57898 237062 58134
rect 237146 57898 237382 58134
rect 236826 22218 237062 22454
rect 237146 22218 237382 22454
rect 236826 21898 237062 22134
rect 237146 21898 237382 22134
rect 236826 -5382 237062 -5146
rect 237146 -5382 237382 -5146
rect 236826 -5702 237062 -5466
rect 237146 -5702 237382 -5466
rect 240546 710362 240782 710598
rect 240866 710362 241102 710598
rect 240546 710042 240782 710278
rect 240866 710042 241102 710278
rect 240546 673938 240782 674174
rect 240866 673938 241102 674174
rect 240546 673618 240782 673854
rect 240866 673618 241102 673854
rect 240546 637938 240782 638174
rect 240866 637938 241102 638174
rect 240546 637618 240782 637854
rect 240866 637618 241102 637854
rect 240546 601938 240782 602174
rect 240866 601938 241102 602174
rect 240546 601618 240782 601854
rect 240866 601618 241102 601854
rect 240546 565938 240782 566174
rect 240866 565938 241102 566174
rect 240546 565618 240782 565854
rect 240866 565618 241102 565854
rect 240546 529938 240782 530174
rect 240866 529938 241102 530174
rect 240546 529618 240782 529854
rect 240866 529618 241102 529854
rect 240546 493938 240782 494174
rect 240866 493938 241102 494174
rect 240546 493618 240782 493854
rect 240866 493618 241102 493854
rect 240546 457938 240782 458174
rect 240866 457938 241102 458174
rect 240546 457618 240782 457854
rect 240866 457618 241102 457854
rect 240546 421938 240782 422174
rect 240866 421938 241102 422174
rect 240546 421618 240782 421854
rect 240866 421618 241102 421854
rect 240546 385938 240782 386174
rect 240866 385938 241102 386174
rect 240546 385618 240782 385854
rect 240866 385618 241102 385854
rect 240546 349938 240782 350174
rect 240866 349938 241102 350174
rect 240546 349618 240782 349854
rect 240866 349618 241102 349854
rect 240546 313938 240782 314174
rect 240866 313938 241102 314174
rect 240546 313618 240782 313854
rect 240866 313618 241102 313854
rect 240546 277938 240782 278174
rect 240866 277938 241102 278174
rect 240546 277618 240782 277854
rect 240866 277618 241102 277854
rect 240546 241938 240782 242174
rect 240866 241938 241102 242174
rect 240546 241618 240782 241854
rect 240866 241618 241102 241854
rect 240546 205938 240782 206174
rect 240866 205938 241102 206174
rect 240546 205618 240782 205854
rect 240866 205618 241102 205854
rect 240546 169938 240782 170174
rect 240866 169938 241102 170174
rect 240546 169618 240782 169854
rect 240866 169618 241102 169854
rect 240546 133938 240782 134174
rect 240866 133938 241102 134174
rect 240546 133618 240782 133854
rect 240866 133618 241102 133854
rect 240546 97938 240782 98174
rect 240866 97938 241102 98174
rect 240546 97618 240782 97854
rect 240866 97618 241102 97854
rect 240546 61938 240782 62174
rect 240866 61938 241102 62174
rect 240546 61618 240782 61854
rect 240866 61618 241102 61854
rect 240546 25938 240782 26174
rect 240866 25938 241102 26174
rect 240546 25618 240782 25854
rect 240866 25618 241102 25854
rect 244266 711322 244502 711558
rect 244586 711322 244822 711558
rect 244266 711002 244502 711238
rect 244586 711002 244822 711238
rect 244266 677658 244502 677894
rect 244586 677658 244822 677894
rect 244266 677338 244502 677574
rect 244586 677338 244822 677574
rect 244266 641658 244502 641894
rect 244586 641658 244822 641894
rect 244266 641338 244502 641574
rect 244586 641338 244822 641574
rect 244266 605658 244502 605894
rect 244586 605658 244822 605894
rect 244266 605338 244502 605574
rect 244586 605338 244822 605574
rect 244266 569658 244502 569894
rect 244586 569658 244822 569894
rect 244266 569338 244502 569574
rect 244586 569338 244822 569574
rect 244266 533658 244502 533894
rect 244586 533658 244822 533894
rect 244266 533338 244502 533574
rect 244586 533338 244822 533574
rect 244266 497658 244502 497894
rect 244586 497658 244822 497894
rect 244266 497338 244502 497574
rect 244586 497338 244822 497574
rect 244266 461658 244502 461894
rect 244586 461658 244822 461894
rect 244266 461338 244502 461574
rect 244586 461338 244822 461574
rect 244266 425658 244502 425894
rect 244586 425658 244822 425894
rect 244266 425338 244502 425574
rect 244586 425338 244822 425574
rect 244266 389658 244502 389894
rect 244586 389658 244822 389894
rect 244266 389338 244502 389574
rect 244586 389338 244822 389574
rect 244266 353658 244502 353894
rect 244586 353658 244822 353894
rect 244266 353338 244502 353574
rect 244586 353338 244822 353574
rect 244266 317658 244502 317894
rect 244586 317658 244822 317894
rect 244266 317338 244502 317574
rect 244586 317338 244822 317574
rect 244266 281658 244502 281894
rect 244586 281658 244822 281894
rect 244266 281338 244502 281574
rect 244586 281338 244822 281574
rect 244266 245658 244502 245894
rect 244586 245658 244822 245894
rect 244266 245338 244502 245574
rect 244586 245338 244822 245574
rect 244266 209658 244502 209894
rect 244586 209658 244822 209894
rect 244266 209338 244502 209574
rect 244586 209338 244822 209574
rect 244266 173658 244502 173894
rect 244586 173658 244822 173894
rect 244266 173338 244502 173574
rect 244586 173338 244822 173574
rect 244266 137658 244502 137894
rect 244586 137658 244822 137894
rect 244266 137338 244502 137574
rect 244586 137338 244822 137574
rect 244266 101658 244502 101894
rect 244586 101658 244822 101894
rect 244266 101338 244502 101574
rect 244586 101338 244822 101574
rect 244266 65658 244502 65894
rect 244586 65658 244822 65894
rect 244266 65338 244502 65574
rect 244586 65338 244822 65574
rect 244266 29658 244502 29894
rect 244586 29658 244822 29894
rect 244266 29338 244502 29574
rect 244586 29338 244822 29574
rect 240546 -6342 240782 -6106
rect 240866 -6342 241102 -6106
rect 240546 -6662 240782 -6426
rect 240866 -6662 241102 -6426
rect 244266 -7302 244502 -7066
rect 244586 -7302 244822 -7066
rect 244266 -7622 244502 -7386
rect 244586 -7622 244822 -7386
rect 254226 704602 254462 704838
rect 254546 704602 254782 704838
rect 254226 704282 254462 704518
rect 254546 704282 254782 704518
rect 254226 687618 254462 687854
rect 254546 687618 254782 687854
rect 254226 687298 254462 687534
rect 254546 687298 254782 687534
rect 254226 651618 254462 651854
rect 254546 651618 254782 651854
rect 254226 651298 254462 651534
rect 254546 651298 254782 651534
rect 254226 615618 254462 615854
rect 254546 615618 254782 615854
rect 254226 615298 254462 615534
rect 254546 615298 254782 615534
rect 254226 579618 254462 579854
rect 254546 579618 254782 579854
rect 254226 579298 254462 579534
rect 254546 579298 254782 579534
rect 254226 543618 254462 543854
rect 254546 543618 254782 543854
rect 254226 543298 254462 543534
rect 254546 543298 254782 543534
rect 254226 507618 254462 507854
rect 254546 507618 254782 507854
rect 254226 507298 254462 507534
rect 254546 507298 254782 507534
rect 254226 471618 254462 471854
rect 254546 471618 254782 471854
rect 254226 471298 254462 471534
rect 254546 471298 254782 471534
rect 254226 435618 254462 435854
rect 254546 435618 254782 435854
rect 254226 435298 254462 435534
rect 254546 435298 254782 435534
rect 254226 399618 254462 399854
rect 254546 399618 254782 399854
rect 254226 399298 254462 399534
rect 254546 399298 254782 399534
rect 254226 363618 254462 363854
rect 254546 363618 254782 363854
rect 254226 363298 254462 363534
rect 254546 363298 254782 363534
rect 254226 327618 254462 327854
rect 254546 327618 254782 327854
rect 254226 327298 254462 327534
rect 254546 327298 254782 327534
rect 254226 291618 254462 291854
rect 254546 291618 254782 291854
rect 254226 291298 254462 291534
rect 254546 291298 254782 291534
rect 254226 255618 254462 255854
rect 254546 255618 254782 255854
rect 254226 255298 254462 255534
rect 254546 255298 254782 255534
rect 254226 219618 254462 219854
rect 254546 219618 254782 219854
rect 254226 219298 254462 219534
rect 254546 219298 254782 219534
rect 254226 183618 254462 183854
rect 254546 183618 254782 183854
rect 254226 183298 254462 183534
rect 254546 183298 254782 183534
rect 254226 147618 254462 147854
rect 254546 147618 254782 147854
rect 254226 147298 254462 147534
rect 254546 147298 254782 147534
rect 254226 111618 254462 111854
rect 254546 111618 254782 111854
rect 254226 111298 254462 111534
rect 254546 111298 254782 111534
rect 254226 75618 254462 75854
rect 254546 75618 254782 75854
rect 254226 75298 254462 75534
rect 254546 75298 254782 75534
rect 254226 39618 254462 39854
rect 254546 39618 254782 39854
rect 254226 39298 254462 39534
rect 254546 39298 254782 39534
rect 254226 3618 254462 3854
rect 254546 3618 254782 3854
rect 254226 3298 254462 3534
rect 254546 3298 254782 3534
rect 254226 -582 254462 -346
rect 254546 -582 254782 -346
rect 254226 -902 254462 -666
rect 254546 -902 254782 -666
rect 257946 705562 258182 705798
rect 258266 705562 258502 705798
rect 257946 705242 258182 705478
rect 258266 705242 258502 705478
rect 257946 691338 258182 691574
rect 258266 691338 258502 691574
rect 257946 691018 258182 691254
rect 258266 691018 258502 691254
rect 257946 655338 258182 655574
rect 258266 655338 258502 655574
rect 257946 655018 258182 655254
rect 258266 655018 258502 655254
rect 257946 619338 258182 619574
rect 258266 619338 258502 619574
rect 257946 619018 258182 619254
rect 258266 619018 258502 619254
rect 257946 583338 258182 583574
rect 258266 583338 258502 583574
rect 257946 583018 258182 583254
rect 258266 583018 258502 583254
rect 257946 547338 258182 547574
rect 258266 547338 258502 547574
rect 257946 547018 258182 547254
rect 258266 547018 258502 547254
rect 257946 511338 258182 511574
rect 258266 511338 258502 511574
rect 257946 511018 258182 511254
rect 258266 511018 258502 511254
rect 257946 475338 258182 475574
rect 258266 475338 258502 475574
rect 257946 475018 258182 475254
rect 258266 475018 258502 475254
rect 257946 439338 258182 439574
rect 258266 439338 258502 439574
rect 257946 439018 258182 439254
rect 258266 439018 258502 439254
rect 257946 403338 258182 403574
rect 258266 403338 258502 403574
rect 257946 403018 258182 403254
rect 258266 403018 258502 403254
rect 257946 367338 258182 367574
rect 258266 367338 258502 367574
rect 257946 367018 258182 367254
rect 258266 367018 258502 367254
rect 257946 331338 258182 331574
rect 258266 331338 258502 331574
rect 257946 331018 258182 331254
rect 258266 331018 258502 331254
rect 257946 295338 258182 295574
rect 258266 295338 258502 295574
rect 257946 295018 258182 295254
rect 258266 295018 258502 295254
rect 257946 259338 258182 259574
rect 258266 259338 258502 259574
rect 257946 259018 258182 259254
rect 258266 259018 258502 259254
rect 257946 223338 258182 223574
rect 258266 223338 258502 223574
rect 257946 223018 258182 223254
rect 258266 223018 258502 223254
rect 257946 187338 258182 187574
rect 258266 187338 258502 187574
rect 257946 187018 258182 187254
rect 258266 187018 258502 187254
rect 257946 151338 258182 151574
rect 258266 151338 258502 151574
rect 257946 151018 258182 151254
rect 258266 151018 258502 151254
rect 257946 115338 258182 115574
rect 258266 115338 258502 115574
rect 257946 115018 258182 115254
rect 258266 115018 258502 115254
rect 257946 79338 258182 79574
rect 258266 79338 258502 79574
rect 257946 79018 258182 79254
rect 258266 79018 258502 79254
rect 257946 43338 258182 43574
rect 258266 43338 258502 43574
rect 257946 43018 258182 43254
rect 258266 43018 258502 43254
rect 257946 7338 258182 7574
rect 258266 7338 258502 7574
rect 257946 7018 258182 7254
rect 258266 7018 258502 7254
rect 257946 -1542 258182 -1306
rect 258266 -1542 258502 -1306
rect 257946 -1862 258182 -1626
rect 258266 -1862 258502 -1626
rect 261666 706522 261902 706758
rect 261986 706522 262222 706758
rect 261666 706202 261902 706438
rect 261986 706202 262222 706438
rect 261666 695058 261902 695294
rect 261986 695058 262222 695294
rect 261666 694738 261902 694974
rect 261986 694738 262222 694974
rect 261666 659058 261902 659294
rect 261986 659058 262222 659294
rect 261666 658738 261902 658974
rect 261986 658738 262222 658974
rect 261666 623058 261902 623294
rect 261986 623058 262222 623294
rect 261666 622738 261902 622974
rect 261986 622738 262222 622974
rect 261666 587058 261902 587294
rect 261986 587058 262222 587294
rect 261666 586738 261902 586974
rect 261986 586738 262222 586974
rect 261666 551058 261902 551294
rect 261986 551058 262222 551294
rect 261666 550738 261902 550974
rect 261986 550738 262222 550974
rect 261666 515058 261902 515294
rect 261986 515058 262222 515294
rect 261666 514738 261902 514974
rect 261986 514738 262222 514974
rect 261666 479058 261902 479294
rect 261986 479058 262222 479294
rect 261666 478738 261902 478974
rect 261986 478738 262222 478974
rect 261666 443058 261902 443294
rect 261986 443058 262222 443294
rect 261666 442738 261902 442974
rect 261986 442738 262222 442974
rect 261666 407058 261902 407294
rect 261986 407058 262222 407294
rect 261666 406738 261902 406974
rect 261986 406738 262222 406974
rect 261666 371058 261902 371294
rect 261986 371058 262222 371294
rect 261666 370738 261902 370974
rect 261986 370738 262222 370974
rect 261666 335058 261902 335294
rect 261986 335058 262222 335294
rect 261666 334738 261902 334974
rect 261986 334738 262222 334974
rect 261666 299058 261902 299294
rect 261986 299058 262222 299294
rect 261666 298738 261902 298974
rect 261986 298738 262222 298974
rect 261666 263058 261902 263294
rect 261986 263058 262222 263294
rect 261666 262738 261902 262974
rect 261986 262738 262222 262974
rect 261666 227058 261902 227294
rect 261986 227058 262222 227294
rect 261666 226738 261902 226974
rect 261986 226738 262222 226974
rect 261666 191058 261902 191294
rect 261986 191058 262222 191294
rect 261666 190738 261902 190974
rect 261986 190738 262222 190974
rect 261666 155058 261902 155294
rect 261986 155058 262222 155294
rect 261666 154738 261902 154974
rect 261986 154738 262222 154974
rect 261666 119058 261902 119294
rect 261986 119058 262222 119294
rect 261666 118738 261902 118974
rect 261986 118738 262222 118974
rect 261666 83058 261902 83294
rect 261986 83058 262222 83294
rect 261666 82738 261902 82974
rect 261986 82738 262222 82974
rect 261666 47058 261902 47294
rect 261986 47058 262222 47294
rect 261666 46738 261902 46974
rect 261986 46738 262222 46974
rect 261666 11058 261902 11294
rect 261986 11058 262222 11294
rect 261666 10738 261902 10974
rect 261986 10738 262222 10974
rect 261666 -2502 261902 -2266
rect 261986 -2502 262222 -2266
rect 261666 -2822 261902 -2586
rect 261986 -2822 262222 -2586
rect 265386 707482 265622 707718
rect 265706 707482 265942 707718
rect 265386 707162 265622 707398
rect 265706 707162 265942 707398
rect 265386 698778 265622 699014
rect 265706 698778 265942 699014
rect 265386 698458 265622 698694
rect 265706 698458 265942 698694
rect 265386 662778 265622 663014
rect 265706 662778 265942 663014
rect 265386 662458 265622 662694
rect 265706 662458 265942 662694
rect 265386 626778 265622 627014
rect 265706 626778 265942 627014
rect 265386 626458 265622 626694
rect 265706 626458 265942 626694
rect 265386 590778 265622 591014
rect 265706 590778 265942 591014
rect 265386 590458 265622 590694
rect 265706 590458 265942 590694
rect 265386 554778 265622 555014
rect 265706 554778 265942 555014
rect 265386 554458 265622 554694
rect 265706 554458 265942 554694
rect 265386 518778 265622 519014
rect 265706 518778 265942 519014
rect 265386 518458 265622 518694
rect 265706 518458 265942 518694
rect 265386 482778 265622 483014
rect 265706 482778 265942 483014
rect 265386 482458 265622 482694
rect 265706 482458 265942 482694
rect 265386 446778 265622 447014
rect 265706 446778 265942 447014
rect 265386 446458 265622 446694
rect 265706 446458 265942 446694
rect 265386 410778 265622 411014
rect 265706 410778 265942 411014
rect 265386 410458 265622 410694
rect 265706 410458 265942 410694
rect 265386 374778 265622 375014
rect 265706 374778 265942 375014
rect 265386 374458 265622 374694
rect 265706 374458 265942 374694
rect 265386 338778 265622 339014
rect 265706 338778 265942 339014
rect 265386 338458 265622 338694
rect 265706 338458 265942 338694
rect 265386 302778 265622 303014
rect 265706 302778 265942 303014
rect 265386 302458 265622 302694
rect 265706 302458 265942 302694
rect 265386 266778 265622 267014
rect 265706 266778 265942 267014
rect 265386 266458 265622 266694
rect 265706 266458 265942 266694
rect 265386 230778 265622 231014
rect 265706 230778 265942 231014
rect 265386 230458 265622 230694
rect 265706 230458 265942 230694
rect 265386 194778 265622 195014
rect 265706 194778 265942 195014
rect 265386 194458 265622 194694
rect 265706 194458 265942 194694
rect 265386 158778 265622 159014
rect 265706 158778 265942 159014
rect 265386 158458 265622 158694
rect 265706 158458 265942 158694
rect 265386 122778 265622 123014
rect 265706 122778 265942 123014
rect 265386 122458 265622 122694
rect 265706 122458 265942 122694
rect 265386 86778 265622 87014
rect 265706 86778 265942 87014
rect 265386 86458 265622 86694
rect 265706 86458 265942 86694
rect 265386 50778 265622 51014
rect 265706 50778 265942 51014
rect 265386 50458 265622 50694
rect 265706 50458 265942 50694
rect 265386 14778 265622 15014
rect 265706 14778 265942 15014
rect 265386 14458 265622 14694
rect 265706 14458 265942 14694
rect 265386 -3462 265622 -3226
rect 265706 -3462 265942 -3226
rect 265386 -3782 265622 -3546
rect 265706 -3782 265942 -3546
rect 269106 708442 269342 708678
rect 269426 708442 269662 708678
rect 269106 708122 269342 708358
rect 269426 708122 269662 708358
rect 269106 666498 269342 666734
rect 269426 666498 269662 666734
rect 269106 666178 269342 666414
rect 269426 666178 269662 666414
rect 269106 630498 269342 630734
rect 269426 630498 269662 630734
rect 269106 630178 269342 630414
rect 269426 630178 269662 630414
rect 269106 594498 269342 594734
rect 269426 594498 269662 594734
rect 269106 594178 269342 594414
rect 269426 594178 269662 594414
rect 269106 558498 269342 558734
rect 269426 558498 269662 558734
rect 269106 558178 269342 558414
rect 269426 558178 269662 558414
rect 269106 522498 269342 522734
rect 269426 522498 269662 522734
rect 269106 522178 269342 522414
rect 269426 522178 269662 522414
rect 269106 486498 269342 486734
rect 269426 486498 269662 486734
rect 269106 486178 269342 486414
rect 269426 486178 269662 486414
rect 269106 450498 269342 450734
rect 269426 450498 269662 450734
rect 269106 450178 269342 450414
rect 269426 450178 269662 450414
rect 269106 414498 269342 414734
rect 269426 414498 269662 414734
rect 269106 414178 269342 414414
rect 269426 414178 269662 414414
rect 269106 378498 269342 378734
rect 269426 378498 269662 378734
rect 269106 378178 269342 378414
rect 269426 378178 269662 378414
rect 269106 342498 269342 342734
rect 269426 342498 269662 342734
rect 269106 342178 269342 342414
rect 269426 342178 269662 342414
rect 269106 306498 269342 306734
rect 269426 306498 269662 306734
rect 269106 306178 269342 306414
rect 269426 306178 269662 306414
rect 269106 270498 269342 270734
rect 269426 270498 269662 270734
rect 269106 270178 269342 270414
rect 269426 270178 269662 270414
rect 269106 234498 269342 234734
rect 269426 234498 269662 234734
rect 269106 234178 269342 234414
rect 269426 234178 269662 234414
rect 269106 198498 269342 198734
rect 269426 198498 269662 198734
rect 269106 198178 269342 198414
rect 269426 198178 269662 198414
rect 269106 162498 269342 162734
rect 269426 162498 269662 162734
rect 269106 162178 269342 162414
rect 269426 162178 269662 162414
rect 269106 126498 269342 126734
rect 269426 126498 269662 126734
rect 269106 126178 269342 126414
rect 269426 126178 269662 126414
rect 269106 90498 269342 90734
rect 269426 90498 269662 90734
rect 269106 90178 269342 90414
rect 269426 90178 269662 90414
rect 269106 54498 269342 54734
rect 269426 54498 269662 54734
rect 269106 54178 269342 54414
rect 269426 54178 269662 54414
rect 269106 18498 269342 18734
rect 269426 18498 269662 18734
rect 269106 18178 269342 18414
rect 269426 18178 269662 18414
rect 269106 -4422 269342 -4186
rect 269426 -4422 269662 -4186
rect 269106 -4742 269342 -4506
rect 269426 -4742 269662 -4506
rect 272826 709402 273062 709638
rect 273146 709402 273382 709638
rect 272826 709082 273062 709318
rect 273146 709082 273382 709318
rect 272826 670218 273062 670454
rect 273146 670218 273382 670454
rect 272826 669898 273062 670134
rect 273146 669898 273382 670134
rect 272826 634218 273062 634454
rect 273146 634218 273382 634454
rect 272826 633898 273062 634134
rect 273146 633898 273382 634134
rect 272826 598218 273062 598454
rect 273146 598218 273382 598454
rect 272826 597898 273062 598134
rect 273146 597898 273382 598134
rect 272826 562218 273062 562454
rect 273146 562218 273382 562454
rect 272826 561898 273062 562134
rect 273146 561898 273382 562134
rect 272826 526218 273062 526454
rect 273146 526218 273382 526454
rect 272826 525898 273062 526134
rect 273146 525898 273382 526134
rect 272826 490218 273062 490454
rect 273146 490218 273382 490454
rect 272826 489898 273062 490134
rect 273146 489898 273382 490134
rect 272826 454218 273062 454454
rect 273146 454218 273382 454454
rect 272826 453898 273062 454134
rect 273146 453898 273382 454134
rect 272826 418218 273062 418454
rect 273146 418218 273382 418454
rect 272826 417898 273062 418134
rect 273146 417898 273382 418134
rect 272826 382218 273062 382454
rect 273146 382218 273382 382454
rect 272826 381898 273062 382134
rect 273146 381898 273382 382134
rect 272826 346218 273062 346454
rect 273146 346218 273382 346454
rect 272826 345898 273062 346134
rect 273146 345898 273382 346134
rect 272826 310218 273062 310454
rect 273146 310218 273382 310454
rect 272826 309898 273062 310134
rect 273146 309898 273382 310134
rect 272826 274218 273062 274454
rect 273146 274218 273382 274454
rect 272826 273898 273062 274134
rect 273146 273898 273382 274134
rect 272826 238218 273062 238454
rect 273146 238218 273382 238454
rect 272826 237898 273062 238134
rect 273146 237898 273382 238134
rect 272826 202218 273062 202454
rect 273146 202218 273382 202454
rect 272826 201898 273062 202134
rect 273146 201898 273382 202134
rect 272826 166218 273062 166454
rect 273146 166218 273382 166454
rect 272826 165898 273062 166134
rect 273146 165898 273382 166134
rect 272826 130218 273062 130454
rect 273146 130218 273382 130454
rect 272826 129898 273062 130134
rect 273146 129898 273382 130134
rect 272826 94218 273062 94454
rect 273146 94218 273382 94454
rect 272826 93898 273062 94134
rect 273146 93898 273382 94134
rect 272826 58218 273062 58454
rect 273146 58218 273382 58454
rect 272826 57898 273062 58134
rect 273146 57898 273382 58134
rect 272826 22218 273062 22454
rect 273146 22218 273382 22454
rect 272826 21898 273062 22134
rect 273146 21898 273382 22134
rect 272826 -5382 273062 -5146
rect 273146 -5382 273382 -5146
rect 272826 -5702 273062 -5466
rect 273146 -5702 273382 -5466
rect 276546 710362 276782 710598
rect 276866 710362 277102 710598
rect 276546 710042 276782 710278
rect 276866 710042 277102 710278
rect 276546 673938 276782 674174
rect 276866 673938 277102 674174
rect 276546 673618 276782 673854
rect 276866 673618 277102 673854
rect 276546 637938 276782 638174
rect 276866 637938 277102 638174
rect 276546 637618 276782 637854
rect 276866 637618 277102 637854
rect 276546 601938 276782 602174
rect 276866 601938 277102 602174
rect 276546 601618 276782 601854
rect 276866 601618 277102 601854
rect 276546 565938 276782 566174
rect 276866 565938 277102 566174
rect 276546 565618 276782 565854
rect 276866 565618 277102 565854
rect 276546 529938 276782 530174
rect 276866 529938 277102 530174
rect 276546 529618 276782 529854
rect 276866 529618 277102 529854
rect 276546 493938 276782 494174
rect 276866 493938 277102 494174
rect 276546 493618 276782 493854
rect 276866 493618 277102 493854
rect 276546 457938 276782 458174
rect 276866 457938 277102 458174
rect 276546 457618 276782 457854
rect 276866 457618 277102 457854
rect 276546 421938 276782 422174
rect 276866 421938 277102 422174
rect 276546 421618 276782 421854
rect 276866 421618 277102 421854
rect 276546 385938 276782 386174
rect 276866 385938 277102 386174
rect 276546 385618 276782 385854
rect 276866 385618 277102 385854
rect 276546 349938 276782 350174
rect 276866 349938 277102 350174
rect 276546 349618 276782 349854
rect 276866 349618 277102 349854
rect 276546 313938 276782 314174
rect 276866 313938 277102 314174
rect 276546 313618 276782 313854
rect 276866 313618 277102 313854
rect 276546 277938 276782 278174
rect 276866 277938 277102 278174
rect 276546 277618 276782 277854
rect 276866 277618 277102 277854
rect 276546 241938 276782 242174
rect 276866 241938 277102 242174
rect 276546 241618 276782 241854
rect 276866 241618 277102 241854
rect 276546 205938 276782 206174
rect 276866 205938 277102 206174
rect 276546 205618 276782 205854
rect 276866 205618 277102 205854
rect 276546 169938 276782 170174
rect 276866 169938 277102 170174
rect 276546 169618 276782 169854
rect 276866 169618 277102 169854
rect 276546 133938 276782 134174
rect 276866 133938 277102 134174
rect 276546 133618 276782 133854
rect 276866 133618 277102 133854
rect 276546 97938 276782 98174
rect 276866 97938 277102 98174
rect 276546 97618 276782 97854
rect 276866 97618 277102 97854
rect 276546 61938 276782 62174
rect 276866 61938 277102 62174
rect 276546 61618 276782 61854
rect 276866 61618 277102 61854
rect 276546 25938 276782 26174
rect 276866 25938 277102 26174
rect 276546 25618 276782 25854
rect 276866 25618 277102 25854
rect 276546 -6342 276782 -6106
rect 276866 -6342 277102 -6106
rect 276546 -6662 276782 -6426
rect 276866 -6662 277102 -6426
rect 280266 711322 280502 711558
rect 280586 711322 280822 711558
rect 280266 711002 280502 711238
rect 280586 711002 280822 711238
rect 280266 677658 280502 677894
rect 280586 677658 280822 677894
rect 280266 677338 280502 677574
rect 280586 677338 280822 677574
rect 280266 641658 280502 641894
rect 280586 641658 280822 641894
rect 280266 641338 280502 641574
rect 280586 641338 280822 641574
rect 280266 605658 280502 605894
rect 280586 605658 280822 605894
rect 280266 605338 280502 605574
rect 280586 605338 280822 605574
rect 280266 569658 280502 569894
rect 280586 569658 280822 569894
rect 280266 569338 280502 569574
rect 280586 569338 280822 569574
rect 280266 533658 280502 533894
rect 280586 533658 280822 533894
rect 280266 533338 280502 533574
rect 280586 533338 280822 533574
rect 280266 497658 280502 497894
rect 280586 497658 280822 497894
rect 280266 497338 280502 497574
rect 280586 497338 280822 497574
rect 280266 461658 280502 461894
rect 280586 461658 280822 461894
rect 280266 461338 280502 461574
rect 280586 461338 280822 461574
rect 280266 425658 280502 425894
rect 280586 425658 280822 425894
rect 280266 425338 280502 425574
rect 280586 425338 280822 425574
rect 280266 389658 280502 389894
rect 280586 389658 280822 389894
rect 280266 389338 280502 389574
rect 280586 389338 280822 389574
rect 280266 353658 280502 353894
rect 280586 353658 280822 353894
rect 280266 353338 280502 353574
rect 280586 353338 280822 353574
rect 280266 317658 280502 317894
rect 280586 317658 280822 317894
rect 280266 317338 280502 317574
rect 280586 317338 280822 317574
rect 280266 281658 280502 281894
rect 280586 281658 280822 281894
rect 280266 281338 280502 281574
rect 280586 281338 280822 281574
rect 280266 245658 280502 245894
rect 280586 245658 280822 245894
rect 280266 245338 280502 245574
rect 280586 245338 280822 245574
rect 280266 209658 280502 209894
rect 280586 209658 280822 209894
rect 280266 209338 280502 209574
rect 280586 209338 280822 209574
rect 280266 173658 280502 173894
rect 280586 173658 280822 173894
rect 280266 173338 280502 173574
rect 280586 173338 280822 173574
rect 280266 137658 280502 137894
rect 280586 137658 280822 137894
rect 280266 137338 280502 137574
rect 280586 137338 280822 137574
rect 280266 101658 280502 101894
rect 280586 101658 280822 101894
rect 280266 101338 280502 101574
rect 280586 101338 280822 101574
rect 280266 65658 280502 65894
rect 280586 65658 280822 65894
rect 280266 65338 280502 65574
rect 280586 65338 280822 65574
rect 280266 29658 280502 29894
rect 280586 29658 280822 29894
rect 280266 29338 280502 29574
rect 280586 29338 280822 29574
rect 280266 -7302 280502 -7066
rect 280586 -7302 280822 -7066
rect 280266 -7622 280502 -7386
rect 280586 -7622 280822 -7386
rect 290226 704602 290462 704838
rect 290546 704602 290782 704838
rect 290226 704282 290462 704518
rect 290546 704282 290782 704518
rect 290226 687618 290462 687854
rect 290546 687618 290782 687854
rect 290226 687298 290462 687534
rect 290546 687298 290782 687534
rect 290226 651618 290462 651854
rect 290546 651618 290782 651854
rect 290226 651298 290462 651534
rect 290546 651298 290782 651534
rect 290226 615618 290462 615854
rect 290546 615618 290782 615854
rect 290226 615298 290462 615534
rect 290546 615298 290782 615534
rect 290226 579618 290462 579854
rect 290546 579618 290782 579854
rect 290226 579298 290462 579534
rect 290546 579298 290782 579534
rect 290226 543618 290462 543854
rect 290546 543618 290782 543854
rect 290226 543298 290462 543534
rect 290546 543298 290782 543534
rect 290226 507618 290462 507854
rect 290546 507618 290782 507854
rect 290226 507298 290462 507534
rect 290546 507298 290782 507534
rect 290226 471618 290462 471854
rect 290546 471618 290782 471854
rect 290226 471298 290462 471534
rect 290546 471298 290782 471534
rect 290226 435618 290462 435854
rect 290546 435618 290782 435854
rect 290226 435298 290462 435534
rect 290546 435298 290782 435534
rect 290226 399618 290462 399854
rect 290546 399618 290782 399854
rect 290226 399298 290462 399534
rect 290546 399298 290782 399534
rect 290226 363618 290462 363854
rect 290546 363618 290782 363854
rect 290226 363298 290462 363534
rect 290546 363298 290782 363534
rect 290226 327618 290462 327854
rect 290546 327618 290782 327854
rect 290226 327298 290462 327534
rect 290546 327298 290782 327534
rect 290226 291618 290462 291854
rect 290546 291618 290782 291854
rect 290226 291298 290462 291534
rect 290546 291298 290782 291534
rect 290226 255618 290462 255854
rect 290546 255618 290782 255854
rect 290226 255298 290462 255534
rect 290546 255298 290782 255534
rect 290226 219618 290462 219854
rect 290546 219618 290782 219854
rect 290226 219298 290462 219534
rect 290546 219298 290782 219534
rect 290226 183618 290462 183854
rect 290546 183618 290782 183854
rect 290226 183298 290462 183534
rect 290546 183298 290782 183534
rect 290226 147618 290462 147854
rect 290546 147618 290782 147854
rect 290226 147298 290462 147534
rect 290546 147298 290782 147534
rect 290226 111618 290462 111854
rect 290546 111618 290782 111854
rect 290226 111298 290462 111534
rect 290546 111298 290782 111534
rect 290226 75618 290462 75854
rect 290546 75618 290782 75854
rect 290226 75298 290462 75534
rect 290546 75298 290782 75534
rect 290226 39618 290462 39854
rect 290546 39618 290782 39854
rect 290226 39298 290462 39534
rect 290546 39298 290782 39534
rect 290226 3618 290462 3854
rect 290546 3618 290782 3854
rect 290226 3298 290462 3534
rect 290546 3298 290782 3534
rect 290226 -582 290462 -346
rect 290546 -582 290782 -346
rect 290226 -902 290462 -666
rect 290546 -902 290782 -666
rect 293946 705562 294182 705798
rect 294266 705562 294502 705798
rect 293946 705242 294182 705478
rect 294266 705242 294502 705478
rect 293946 691338 294182 691574
rect 294266 691338 294502 691574
rect 293946 691018 294182 691254
rect 294266 691018 294502 691254
rect 293946 655338 294182 655574
rect 294266 655338 294502 655574
rect 293946 655018 294182 655254
rect 294266 655018 294502 655254
rect 293946 619338 294182 619574
rect 294266 619338 294502 619574
rect 293946 619018 294182 619254
rect 294266 619018 294502 619254
rect 293946 583338 294182 583574
rect 294266 583338 294502 583574
rect 293946 583018 294182 583254
rect 294266 583018 294502 583254
rect 293946 547338 294182 547574
rect 294266 547338 294502 547574
rect 293946 547018 294182 547254
rect 294266 547018 294502 547254
rect 293946 511338 294182 511574
rect 294266 511338 294502 511574
rect 293946 511018 294182 511254
rect 294266 511018 294502 511254
rect 293946 475338 294182 475574
rect 294266 475338 294502 475574
rect 293946 475018 294182 475254
rect 294266 475018 294502 475254
rect 293946 439338 294182 439574
rect 294266 439338 294502 439574
rect 293946 439018 294182 439254
rect 294266 439018 294502 439254
rect 293946 403338 294182 403574
rect 294266 403338 294502 403574
rect 293946 403018 294182 403254
rect 294266 403018 294502 403254
rect 293946 367338 294182 367574
rect 294266 367338 294502 367574
rect 293946 367018 294182 367254
rect 294266 367018 294502 367254
rect 293946 331338 294182 331574
rect 294266 331338 294502 331574
rect 293946 331018 294182 331254
rect 294266 331018 294502 331254
rect 293946 295338 294182 295574
rect 294266 295338 294502 295574
rect 293946 295018 294182 295254
rect 294266 295018 294502 295254
rect 293946 259338 294182 259574
rect 294266 259338 294502 259574
rect 293946 259018 294182 259254
rect 294266 259018 294502 259254
rect 293946 223338 294182 223574
rect 294266 223338 294502 223574
rect 293946 223018 294182 223254
rect 294266 223018 294502 223254
rect 293946 187338 294182 187574
rect 294266 187338 294502 187574
rect 293946 187018 294182 187254
rect 294266 187018 294502 187254
rect 293946 151338 294182 151574
rect 294266 151338 294502 151574
rect 293946 151018 294182 151254
rect 294266 151018 294502 151254
rect 293946 115338 294182 115574
rect 294266 115338 294502 115574
rect 293946 115018 294182 115254
rect 294266 115018 294502 115254
rect 293946 79338 294182 79574
rect 294266 79338 294502 79574
rect 293946 79018 294182 79254
rect 294266 79018 294502 79254
rect 293946 43338 294182 43574
rect 294266 43338 294502 43574
rect 293946 43018 294182 43254
rect 294266 43018 294502 43254
rect 297666 706522 297902 706758
rect 297986 706522 298222 706758
rect 297666 706202 297902 706438
rect 297986 706202 298222 706438
rect 297666 695058 297902 695294
rect 297986 695058 298222 695294
rect 297666 694738 297902 694974
rect 297986 694738 298222 694974
rect 297666 659058 297902 659294
rect 297986 659058 298222 659294
rect 297666 658738 297902 658974
rect 297986 658738 298222 658974
rect 297666 623058 297902 623294
rect 297986 623058 298222 623294
rect 297666 622738 297902 622974
rect 297986 622738 298222 622974
rect 297666 587058 297902 587294
rect 297986 587058 298222 587294
rect 297666 586738 297902 586974
rect 297986 586738 298222 586974
rect 297666 551058 297902 551294
rect 297986 551058 298222 551294
rect 297666 550738 297902 550974
rect 297986 550738 298222 550974
rect 297666 515058 297902 515294
rect 297986 515058 298222 515294
rect 297666 514738 297902 514974
rect 297986 514738 298222 514974
rect 297666 479058 297902 479294
rect 297986 479058 298222 479294
rect 297666 478738 297902 478974
rect 297986 478738 298222 478974
rect 297666 443058 297902 443294
rect 297986 443058 298222 443294
rect 297666 442738 297902 442974
rect 297986 442738 298222 442974
rect 297666 407058 297902 407294
rect 297986 407058 298222 407294
rect 297666 406738 297902 406974
rect 297986 406738 298222 406974
rect 297666 371058 297902 371294
rect 297986 371058 298222 371294
rect 297666 370738 297902 370974
rect 297986 370738 298222 370974
rect 297666 335058 297902 335294
rect 297986 335058 298222 335294
rect 297666 334738 297902 334974
rect 297986 334738 298222 334974
rect 297666 299058 297902 299294
rect 297986 299058 298222 299294
rect 297666 298738 297902 298974
rect 297986 298738 298222 298974
rect 297666 263058 297902 263294
rect 297986 263058 298222 263294
rect 297666 262738 297902 262974
rect 297986 262738 298222 262974
rect 297666 227058 297902 227294
rect 297986 227058 298222 227294
rect 297666 226738 297902 226974
rect 297986 226738 298222 226974
rect 297666 191058 297902 191294
rect 297986 191058 298222 191294
rect 297666 190738 297902 190974
rect 297986 190738 298222 190974
rect 297666 155058 297902 155294
rect 297986 155058 298222 155294
rect 297666 154738 297902 154974
rect 297986 154738 298222 154974
rect 297666 119058 297902 119294
rect 297986 119058 298222 119294
rect 297666 118738 297902 118974
rect 297986 118738 298222 118974
rect 297666 83058 297902 83294
rect 297986 83058 298222 83294
rect 297666 82738 297902 82974
rect 297986 82738 298222 82974
rect 297666 47058 297902 47294
rect 297986 47058 298222 47294
rect 297666 46738 297902 46974
rect 297986 46738 298222 46974
rect 297666 11058 297902 11294
rect 297986 11058 298222 11294
rect 297666 10738 297902 10974
rect 297986 10738 298222 10974
rect 296582 8382 296818 8618
rect 293946 7338 294182 7574
rect 294266 7338 294502 7574
rect 293946 7018 294182 7254
rect 294266 7018 294502 7254
rect 293946 -1542 294182 -1306
rect 294266 -1542 294502 -1306
rect 293946 -1862 294182 -1626
rect 294266 -1862 294502 -1626
rect 297666 -2502 297902 -2266
rect 297986 -2502 298222 -2266
rect 297666 -2822 297902 -2586
rect 297986 -2822 298222 -2586
rect 301386 707482 301622 707718
rect 301706 707482 301942 707718
rect 301386 707162 301622 707398
rect 301706 707162 301942 707398
rect 301386 698778 301622 699014
rect 301706 698778 301942 699014
rect 301386 698458 301622 698694
rect 301706 698458 301942 698694
rect 301386 662778 301622 663014
rect 301706 662778 301942 663014
rect 301386 662458 301622 662694
rect 301706 662458 301942 662694
rect 301386 626778 301622 627014
rect 301706 626778 301942 627014
rect 301386 626458 301622 626694
rect 301706 626458 301942 626694
rect 301386 590778 301622 591014
rect 301706 590778 301942 591014
rect 301386 590458 301622 590694
rect 301706 590458 301942 590694
rect 301386 554778 301622 555014
rect 301706 554778 301942 555014
rect 301386 554458 301622 554694
rect 301706 554458 301942 554694
rect 301386 518778 301622 519014
rect 301706 518778 301942 519014
rect 301386 518458 301622 518694
rect 301706 518458 301942 518694
rect 301386 482778 301622 483014
rect 301706 482778 301942 483014
rect 301386 482458 301622 482694
rect 301706 482458 301942 482694
rect 301386 446778 301622 447014
rect 301706 446778 301942 447014
rect 301386 446458 301622 446694
rect 301706 446458 301942 446694
rect 301386 410778 301622 411014
rect 301706 410778 301942 411014
rect 301386 410458 301622 410694
rect 301706 410458 301942 410694
rect 301386 374778 301622 375014
rect 301706 374778 301942 375014
rect 301386 374458 301622 374694
rect 301706 374458 301942 374694
rect 301386 338778 301622 339014
rect 301706 338778 301942 339014
rect 301386 338458 301622 338694
rect 301706 338458 301942 338694
rect 301386 302778 301622 303014
rect 301706 302778 301942 303014
rect 301386 302458 301622 302694
rect 301706 302458 301942 302694
rect 301386 266778 301622 267014
rect 301706 266778 301942 267014
rect 301386 266458 301622 266694
rect 301706 266458 301942 266694
rect 301386 230778 301622 231014
rect 301706 230778 301942 231014
rect 301386 230458 301622 230694
rect 301706 230458 301942 230694
rect 301386 194778 301622 195014
rect 301706 194778 301942 195014
rect 301386 194458 301622 194694
rect 301706 194458 301942 194694
rect 301386 158778 301622 159014
rect 301706 158778 301942 159014
rect 301386 158458 301622 158694
rect 301706 158458 301942 158694
rect 301386 122778 301622 123014
rect 301706 122778 301942 123014
rect 301386 122458 301622 122694
rect 301706 122458 301942 122694
rect 305106 708442 305342 708678
rect 305426 708442 305662 708678
rect 305106 708122 305342 708358
rect 305426 708122 305662 708358
rect 305106 666498 305342 666734
rect 305426 666498 305662 666734
rect 305106 666178 305342 666414
rect 305426 666178 305662 666414
rect 305106 630498 305342 630734
rect 305426 630498 305662 630734
rect 305106 630178 305342 630414
rect 305426 630178 305662 630414
rect 305106 594498 305342 594734
rect 305426 594498 305662 594734
rect 305106 594178 305342 594414
rect 305426 594178 305662 594414
rect 305106 558498 305342 558734
rect 305426 558498 305662 558734
rect 305106 558178 305342 558414
rect 305426 558178 305662 558414
rect 305106 522498 305342 522734
rect 305426 522498 305662 522734
rect 305106 522178 305342 522414
rect 305426 522178 305662 522414
rect 305106 486498 305342 486734
rect 305426 486498 305662 486734
rect 305106 486178 305342 486414
rect 305426 486178 305662 486414
rect 305106 450498 305342 450734
rect 305426 450498 305662 450734
rect 305106 450178 305342 450414
rect 305426 450178 305662 450414
rect 305106 414498 305342 414734
rect 305426 414498 305662 414734
rect 305106 414178 305342 414414
rect 305426 414178 305662 414414
rect 305106 378498 305342 378734
rect 305426 378498 305662 378734
rect 305106 378178 305342 378414
rect 305426 378178 305662 378414
rect 305106 342498 305342 342734
rect 305426 342498 305662 342734
rect 305106 342178 305342 342414
rect 305426 342178 305662 342414
rect 305106 306498 305342 306734
rect 305426 306498 305662 306734
rect 305106 306178 305342 306414
rect 305426 306178 305662 306414
rect 305106 270498 305342 270734
rect 305426 270498 305662 270734
rect 305106 270178 305342 270414
rect 305426 270178 305662 270414
rect 305106 234498 305342 234734
rect 305426 234498 305662 234734
rect 305106 234178 305342 234414
rect 305426 234178 305662 234414
rect 305106 198498 305342 198734
rect 305426 198498 305662 198734
rect 305106 198178 305342 198414
rect 305426 198178 305662 198414
rect 305106 162498 305342 162734
rect 305426 162498 305662 162734
rect 305106 162178 305342 162414
rect 305426 162178 305662 162414
rect 305106 126498 305342 126734
rect 305426 126498 305662 126734
rect 305106 126178 305342 126414
rect 305426 126178 305662 126414
rect 304250 111618 304486 111854
rect 304250 111298 304486 111534
rect 301386 86778 301622 87014
rect 301706 86778 301942 87014
rect 301386 86458 301622 86694
rect 301706 86458 301942 86694
rect 301386 50778 301622 51014
rect 301706 50778 301942 51014
rect 301386 50458 301622 50694
rect 301706 50458 301942 50694
rect 301386 14778 301622 15014
rect 301706 14778 301942 15014
rect 301386 14458 301622 14694
rect 301706 14458 301942 14694
rect 301386 -3462 301622 -3226
rect 301706 -3462 301942 -3226
rect 301386 -3782 301622 -3546
rect 301706 -3782 301942 -3546
rect 305106 90498 305342 90734
rect 305426 90498 305662 90734
rect 305106 90178 305342 90414
rect 305426 90178 305662 90414
rect 305106 54498 305342 54734
rect 305426 54498 305662 54734
rect 305106 54178 305342 54414
rect 305426 54178 305662 54414
rect 305106 18498 305342 18734
rect 305426 18498 305662 18734
rect 305106 18178 305342 18414
rect 305426 18178 305662 18414
rect 305106 -4422 305342 -4186
rect 305426 -4422 305662 -4186
rect 305106 -4742 305342 -4506
rect 305426 -4742 305662 -4506
rect 308826 709402 309062 709638
rect 309146 709402 309382 709638
rect 308826 709082 309062 709318
rect 309146 709082 309382 709318
rect 308826 670218 309062 670454
rect 309146 670218 309382 670454
rect 308826 669898 309062 670134
rect 309146 669898 309382 670134
rect 308826 634218 309062 634454
rect 309146 634218 309382 634454
rect 308826 633898 309062 634134
rect 309146 633898 309382 634134
rect 308826 598218 309062 598454
rect 309146 598218 309382 598454
rect 308826 597898 309062 598134
rect 309146 597898 309382 598134
rect 308826 562218 309062 562454
rect 309146 562218 309382 562454
rect 308826 561898 309062 562134
rect 309146 561898 309382 562134
rect 308826 526218 309062 526454
rect 309146 526218 309382 526454
rect 308826 525898 309062 526134
rect 309146 525898 309382 526134
rect 308826 490218 309062 490454
rect 309146 490218 309382 490454
rect 308826 489898 309062 490134
rect 309146 489898 309382 490134
rect 308826 454218 309062 454454
rect 309146 454218 309382 454454
rect 308826 453898 309062 454134
rect 309146 453898 309382 454134
rect 308826 418218 309062 418454
rect 309146 418218 309382 418454
rect 308826 417898 309062 418134
rect 309146 417898 309382 418134
rect 308826 382218 309062 382454
rect 309146 382218 309382 382454
rect 308826 381898 309062 382134
rect 309146 381898 309382 382134
rect 308826 346218 309062 346454
rect 309146 346218 309382 346454
rect 308826 345898 309062 346134
rect 309146 345898 309382 346134
rect 308826 310218 309062 310454
rect 309146 310218 309382 310454
rect 308826 309898 309062 310134
rect 309146 309898 309382 310134
rect 308826 274218 309062 274454
rect 309146 274218 309382 274454
rect 308826 273898 309062 274134
rect 309146 273898 309382 274134
rect 308826 238218 309062 238454
rect 309146 238218 309382 238454
rect 308826 237898 309062 238134
rect 309146 237898 309382 238134
rect 308826 202218 309062 202454
rect 309146 202218 309382 202454
rect 308826 201898 309062 202134
rect 309146 201898 309382 202134
rect 308826 166218 309062 166454
rect 309146 166218 309382 166454
rect 308826 165898 309062 166134
rect 309146 165898 309382 166134
rect 308826 130218 309062 130454
rect 309146 130218 309382 130454
rect 308826 129898 309062 130134
rect 309146 129898 309382 130134
rect 308826 94218 309062 94454
rect 309146 94218 309382 94454
rect 308826 93898 309062 94134
rect 309146 93898 309382 94134
rect 308826 58218 309062 58454
rect 309146 58218 309382 58454
rect 308826 57898 309062 58134
rect 309146 57898 309382 58134
rect 308826 22218 309062 22454
rect 309146 22218 309382 22454
rect 308826 21898 309062 22134
rect 309146 21898 309382 22134
rect 308826 -5382 309062 -5146
rect 309146 -5382 309382 -5146
rect 308826 -5702 309062 -5466
rect 309146 -5702 309382 -5466
rect 312546 710362 312782 710598
rect 312866 710362 313102 710598
rect 312546 710042 312782 710278
rect 312866 710042 313102 710278
rect 312546 673938 312782 674174
rect 312866 673938 313102 674174
rect 312546 673618 312782 673854
rect 312866 673618 313102 673854
rect 312546 637938 312782 638174
rect 312866 637938 313102 638174
rect 312546 637618 312782 637854
rect 312866 637618 313102 637854
rect 312546 601938 312782 602174
rect 312866 601938 313102 602174
rect 312546 601618 312782 601854
rect 312866 601618 313102 601854
rect 312546 565938 312782 566174
rect 312866 565938 313102 566174
rect 312546 565618 312782 565854
rect 312866 565618 313102 565854
rect 312546 529938 312782 530174
rect 312866 529938 313102 530174
rect 312546 529618 312782 529854
rect 312866 529618 313102 529854
rect 312546 493938 312782 494174
rect 312866 493938 313102 494174
rect 312546 493618 312782 493854
rect 312866 493618 313102 493854
rect 312546 457938 312782 458174
rect 312866 457938 313102 458174
rect 312546 457618 312782 457854
rect 312866 457618 313102 457854
rect 312546 421938 312782 422174
rect 312866 421938 313102 422174
rect 312546 421618 312782 421854
rect 312866 421618 313102 421854
rect 312546 385938 312782 386174
rect 312866 385938 313102 386174
rect 312546 385618 312782 385854
rect 312866 385618 313102 385854
rect 312546 349938 312782 350174
rect 312866 349938 313102 350174
rect 312546 349618 312782 349854
rect 312866 349618 313102 349854
rect 312546 313938 312782 314174
rect 312866 313938 313102 314174
rect 312546 313618 312782 313854
rect 312866 313618 313102 313854
rect 312546 277938 312782 278174
rect 312866 277938 313102 278174
rect 312546 277618 312782 277854
rect 312866 277618 313102 277854
rect 312546 241938 312782 242174
rect 312866 241938 313102 242174
rect 312546 241618 312782 241854
rect 312866 241618 313102 241854
rect 312546 205938 312782 206174
rect 312866 205938 313102 206174
rect 312546 205618 312782 205854
rect 312866 205618 313102 205854
rect 312546 169938 312782 170174
rect 312866 169938 313102 170174
rect 312546 169618 312782 169854
rect 312866 169618 313102 169854
rect 312546 133938 312782 134174
rect 312866 133938 313102 134174
rect 312546 133618 312782 133854
rect 312866 133618 313102 133854
rect 312546 97938 312782 98174
rect 312866 97938 313102 98174
rect 312546 97618 312782 97854
rect 312866 97618 313102 97854
rect 312546 61938 312782 62174
rect 312866 61938 313102 62174
rect 312546 61618 312782 61854
rect 312866 61618 313102 61854
rect 312546 25938 312782 26174
rect 312866 25938 313102 26174
rect 312546 25618 312782 25854
rect 312866 25618 313102 25854
rect 312546 -6342 312782 -6106
rect 312866 -6342 313102 -6106
rect 312546 -6662 312782 -6426
rect 312866 -6662 313102 -6426
rect 316266 711322 316502 711558
rect 316586 711322 316822 711558
rect 316266 711002 316502 711238
rect 316586 711002 316822 711238
rect 316266 677658 316502 677894
rect 316586 677658 316822 677894
rect 316266 677338 316502 677574
rect 316586 677338 316822 677574
rect 316266 641658 316502 641894
rect 316586 641658 316822 641894
rect 316266 641338 316502 641574
rect 316586 641338 316822 641574
rect 316266 605658 316502 605894
rect 316586 605658 316822 605894
rect 316266 605338 316502 605574
rect 316586 605338 316822 605574
rect 316266 569658 316502 569894
rect 316586 569658 316822 569894
rect 316266 569338 316502 569574
rect 316586 569338 316822 569574
rect 316266 533658 316502 533894
rect 316586 533658 316822 533894
rect 316266 533338 316502 533574
rect 316586 533338 316822 533574
rect 316266 497658 316502 497894
rect 316586 497658 316822 497894
rect 316266 497338 316502 497574
rect 316586 497338 316822 497574
rect 316266 461658 316502 461894
rect 316586 461658 316822 461894
rect 316266 461338 316502 461574
rect 316586 461338 316822 461574
rect 316266 425658 316502 425894
rect 316586 425658 316822 425894
rect 316266 425338 316502 425574
rect 316586 425338 316822 425574
rect 316266 389658 316502 389894
rect 316586 389658 316822 389894
rect 316266 389338 316502 389574
rect 316586 389338 316822 389574
rect 316266 353658 316502 353894
rect 316586 353658 316822 353894
rect 316266 353338 316502 353574
rect 316586 353338 316822 353574
rect 316266 317658 316502 317894
rect 316586 317658 316822 317894
rect 316266 317338 316502 317574
rect 316586 317338 316822 317574
rect 316266 281658 316502 281894
rect 316586 281658 316822 281894
rect 316266 281338 316502 281574
rect 316586 281338 316822 281574
rect 316266 245658 316502 245894
rect 316586 245658 316822 245894
rect 316266 245338 316502 245574
rect 316586 245338 316822 245574
rect 316266 209658 316502 209894
rect 316586 209658 316822 209894
rect 316266 209338 316502 209574
rect 316586 209338 316822 209574
rect 316266 173658 316502 173894
rect 316586 173658 316822 173894
rect 316266 173338 316502 173574
rect 316586 173338 316822 173574
rect 316266 137658 316502 137894
rect 316586 137658 316822 137894
rect 316266 137338 316502 137574
rect 316586 137338 316822 137574
rect 326226 704602 326462 704838
rect 326546 704602 326782 704838
rect 326226 704282 326462 704518
rect 326546 704282 326782 704518
rect 326226 687618 326462 687854
rect 326546 687618 326782 687854
rect 326226 687298 326462 687534
rect 326546 687298 326782 687534
rect 326226 651618 326462 651854
rect 326546 651618 326782 651854
rect 326226 651298 326462 651534
rect 326546 651298 326782 651534
rect 326226 615618 326462 615854
rect 326546 615618 326782 615854
rect 326226 615298 326462 615534
rect 326546 615298 326782 615534
rect 326226 579618 326462 579854
rect 326546 579618 326782 579854
rect 326226 579298 326462 579534
rect 326546 579298 326782 579534
rect 326226 543618 326462 543854
rect 326546 543618 326782 543854
rect 326226 543298 326462 543534
rect 326546 543298 326782 543534
rect 326226 507618 326462 507854
rect 326546 507618 326782 507854
rect 326226 507298 326462 507534
rect 326546 507298 326782 507534
rect 326226 471618 326462 471854
rect 326546 471618 326782 471854
rect 326226 471298 326462 471534
rect 326546 471298 326782 471534
rect 326226 435618 326462 435854
rect 326546 435618 326782 435854
rect 326226 435298 326462 435534
rect 326546 435298 326782 435534
rect 326226 399618 326462 399854
rect 326546 399618 326782 399854
rect 326226 399298 326462 399534
rect 326546 399298 326782 399534
rect 326226 363618 326462 363854
rect 326546 363618 326782 363854
rect 326226 363298 326462 363534
rect 326546 363298 326782 363534
rect 326226 327618 326462 327854
rect 326546 327618 326782 327854
rect 326226 327298 326462 327534
rect 326546 327298 326782 327534
rect 326226 291618 326462 291854
rect 326546 291618 326782 291854
rect 326226 291298 326462 291534
rect 326546 291298 326782 291534
rect 326226 255618 326462 255854
rect 326546 255618 326782 255854
rect 326226 255298 326462 255534
rect 326546 255298 326782 255534
rect 326226 219618 326462 219854
rect 326546 219618 326782 219854
rect 326226 219298 326462 219534
rect 326546 219298 326782 219534
rect 326226 183618 326462 183854
rect 326546 183618 326782 183854
rect 326226 183298 326462 183534
rect 326546 183298 326782 183534
rect 326226 147618 326462 147854
rect 326546 147618 326782 147854
rect 326226 147298 326462 147534
rect 326546 147298 326782 147534
rect 319610 115338 319846 115574
rect 319610 115018 319846 115254
rect 316266 101658 316502 101894
rect 316586 101658 316822 101894
rect 316266 101338 316502 101574
rect 316586 101338 316822 101574
rect 326226 111618 326462 111854
rect 326546 111618 326782 111854
rect 326226 111298 326462 111534
rect 326546 111298 326782 111534
rect 324182 77742 324418 77978
rect 316266 65658 316502 65894
rect 316586 65658 316822 65894
rect 316266 65338 316502 65574
rect 316586 65338 316822 65574
rect 316266 29658 316502 29894
rect 316586 29658 316822 29894
rect 316266 29338 316502 29574
rect 316586 29338 316822 29574
rect 316266 -7302 316502 -7066
rect 316586 -7302 316822 -7066
rect 316266 -7622 316502 -7386
rect 316586 -7622 316822 -7386
rect 326226 75618 326462 75854
rect 326546 75618 326782 75854
rect 326226 75298 326462 75534
rect 326546 75298 326782 75534
rect 326226 39618 326462 39854
rect 326546 39618 326782 39854
rect 326226 39298 326462 39534
rect 326546 39298 326782 39534
rect 326226 3618 326462 3854
rect 326546 3618 326782 3854
rect 326226 3298 326462 3534
rect 326546 3298 326782 3534
rect 326226 -582 326462 -346
rect 326546 -582 326782 -346
rect 326226 -902 326462 -666
rect 326546 -902 326782 -666
rect 329946 705562 330182 705798
rect 330266 705562 330502 705798
rect 329946 705242 330182 705478
rect 330266 705242 330502 705478
rect 329946 691338 330182 691574
rect 330266 691338 330502 691574
rect 329946 691018 330182 691254
rect 330266 691018 330502 691254
rect 329946 655338 330182 655574
rect 330266 655338 330502 655574
rect 329946 655018 330182 655254
rect 330266 655018 330502 655254
rect 329946 619338 330182 619574
rect 330266 619338 330502 619574
rect 329946 619018 330182 619254
rect 330266 619018 330502 619254
rect 329946 583338 330182 583574
rect 330266 583338 330502 583574
rect 329946 583018 330182 583254
rect 330266 583018 330502 583254
rect 329946 547338 330182 547574
rect 330266 547338 330502 547574
rect 329946 547018 330182 547254
rect 330266 547018 330502 547254
rect 329946 511338 330182 511574
rect 330266 511338 330502 511574
rect 329946 511018 330182 511254
rect 330266 511018 330502 511254
rect 329946 475338 330182 475574
rect 330266 475338 330502 475574
rect 329946 475018 330182 475254
rect 330266 475018 330502 475254
rect 329946 439338 330182 439574
rect 330266 439338 330502 439574
rect 329946 439018 330182 439254
rect 330266 439018 330502 439254
rect 329946 403338 330182 403574
rect 330266 403338 330502 403574
rect 329946 403018 330182 403254
rect 330266 403018 330502 403254
rect 329946 367338 330182 367574
rect 330266 367338 330502 367574
rect 329946 367018 330182 367254
rect 330266 367018 330502 367254
rect 329946 331338 330182 331574
rect 330266 331338 330502 331574
rect 329946 331018 330182 331254
rect 330266 331018 330502 331254
rect 329946 295338 330182 295574
rect 330266 295338 330502 295574
rect 329946 295018 330182 295254
rect 330266 295018 330502 295254
rect 329946 259338 330182 259574
rect 330266 259338 330502 259574
rect 329946 259018 330182 259254
rect 330266 259018 330502 259254
rect 329946 223338 330182 223574
rect 330266 223338 330502 223574
rect 329946 223018 330182 223254
rect 330266 223018 330502 223254
rect 329946 187338 330182 187574
rect 330266 187338 330502 187574
rect 329946 187018 330182 187254
rect 330266 187018 330502 187254
rect 329946 151338 330182 151574
rect 330266 151338 330502 151574
rect 329946 151018 330182 151254
rect 330266 151018 330502 151254
rect 329946 115338 330182 115574
rect 330266 115338 330502 115574
rect 329946 115018 330182 115254
rect 330266 115018 330502 115254
rect 329946 79338 330182 79574
rect 330266 79338 330502 79574
rect 329946 79018 330182 79254
rect 330266 79018 330502 79254
rect 329946 43338 330182 43574
rect 330266 43338 330502 43574
rect 329946 43018 330182 43254
rect 330266 43018 330502 43254
rect 329946 7338 330182 7574
rect 330266 7338 330502 7574
rect 329946 7018 330182 7254
rect 330266 7018 330502 7254
rect 329946 -1542 330182 -1306
rect 330266 -1542 330502 -1306
rect 329946 -1862 330182 -1626
rect 330266 -1862 330502 -1626
rect 333666 706522 333902 706758
rect 333986 706522 334222 706758
rect 333666 706202 333902 706438
rect 333986 706202 334222 706438
rect 333666 695058 333902 695294
rect 333986 695058 334222 695294
rect 333666 694738 333902 694974
rect 333986 694738 334222 694974
rect 333666 659058 333902 659294
rect 333986 659058 334222 659294
rect 333666 658738 333902 658974
rect 333986 658738 334222 658974
rect 333666 623058 333902 623294
rect 333986 623058 334222 623294
rect 333666 622738 333902 622974
rect 333986 622738 334222 622974
rect 333666 587058 333902 587294
rect 333986 587058 334222 587294
rect 333666 586738 333902 586974
rect 333986 586738 334222 586974
rect 333666 551058 333902 551294
rect 333986 551058 334222 551294
rect 333666 550738 333902 550974
rect 333986 550738 334222 550974
rect 333666 515058 333902 515294
rect 333986 515058 334222 515294
rect 333666 514738 333902 514974
rect 333986 514738 334222 514974
rect 333666 479058 333902 479294
rect 333986 479058 334222 479294
rect 333666 478738 333902 478974
rect 333986 478738 334222 478974
rect 333666 443058 333902 443294
rect 333986 443058 334222 443294
rect 333666 442738 333902 442974
rect 333986 442738 334222 442974
rect 333666 407058 333902 407294
rect 333986 407058 334222 407294
rect 333666 406738 333902 406974
rect 333986 406738 334222 406974
rect 333666 371058 333902 371294
rect 333986 371058 334222 371294
rect 333666 370738 333902 370974
rect 333986 370738 334222 370974
rect 333666 335058 333902 335294
rect 333986 335058 334222 335294
rect 333666 334738 333902 334974
rect 333986 334738 334222 334974
rect 333666 299058 333902 299294
rect 333986 299058 334222 299294
rect 333666 298738 333902 298974
rect 333986 298738 334222 298974
rect 333666 263058 333902 263294
rect 333986 263058 334222 263294
rect 333666 262738 333902 262974
rect 333986 262738 334222 262974
rect 333666 227058 333902 227294
rect 333986 227058 334222 227294
rect 333666 226738 333902 226974
rect 333986 226738 334222 226974
rect 333666 191058 333902 191294
rect 333986 191058 334222 191294
rect 333666 190738 333902 190974
rect 333986 190738 334222 190974
rect 333666 155058 333902 155294
rect 333986 155058 334222 155294
rect 333666 154738 333902 154974
rect 333986 154738 334222 154974
rect 333666 119058 333902 119294
rect 333986 119058 334222 119294
rect 333666 118738 333902 118974
rect 333986 118738 334222 118974
rect 337386 707482 337622 707718
rect 337706 707482 337942 707718
rect 337386 707162 337622 707398
rect 337706 707162 337942 707398
rect 337386 698778 337622 699014
rect 337706 698778 337942 699014
rect 337386 698458 337622 698694
rect 337706 698458 337942 698694
rect 337386 662778 337622 663014
rect 337706 662778 337942 663014
rect 337386 662458 337622 662694
rect 337706 662458 337942 662694
rect 337386 626778 337622 627014
rect 337706 626778 337942 627014
rect 337386 626458 337622 626694
rect 337706 626458 337942 626694
rect 337386 590778 337622 591014
rect 337706 590778 337942 591014
rect 337386 590458 337622 590694
rect 337706 590458 337942 590694
rect 337386 554778 337622 555014
rect 337706 554778 337942 555014
rect 337386 554458 337622 554694
rect 337706 554458 337942 554694
rect 337386 518778 337622 519014
rect 337706 518778 337942 519014
rect 337386 518458 337622 518694
rect 337706 518458 337942 518694
rect 337386 482778 337622 483014
rect 337706 482778 337942 483014
rect 337386 482458 337622 482694
rect 337706 482458 337942 482694
rect 337386 446778 337622 447014
rect 337706 446778 337942 447014
rect 337386 446458 337622 446694
rect 337706 446458 337942 446694
rect 337386 410778 337622 411014
rect 337706 410778 337942 411014
rect 337386 410458 337622 410694
rect 337706 410458 337942 410694
rect 337386 374778 337622 375014
rect 337706 374778 337942 375014
rect 337386 374458 337622 374694
rect 337706 374458 337942 374694
rect 337386 338778 337622 339014
rect 337706 338778 337942 339014
rect 337386 338458 337622 338694
rect 337706 338458 337942 338694
rect 337386 302778 337622 303014
rect 337706 302778 337942 303014
rect 337386 302458 337622 302694
rect 337706 302458 337942 302694
rect 337386 266778 337622 267014
rect 337706 266778 337942 267014
rect 337386 266458 337622 266694
rect 337706 266458 337942 266694
rect 337386 230778 337622 231014
rect 337706 230778 337942 231014
rect 337386 230458 337622 230694
rect 337706 230458 337942 230694
rect 337386 194778 337622 195014
rect 337706 194778 337942 195014
rect 337386 194458 337622 194694
rect 337706 194458 337942 194694
rect 337386 158778 337622 159014
rect 337706 158778 337942 159014
rect 337386 158458 337622 158694
rect 337706 158458 337942 158694
rect 337386 122778 337622 123014
rect 337706 122778 337942 123014
rect 337386 122458 337622 122694
rect 337706 122458 337942 122694
rect 334970 111618 335206 111854
rect 334970 111298 335206 111534
rect 333666 83058 333902 83294
rect 333986 83058 334222 83294
rect 333666 82738 333902 82974
rect 333986 82738 334222 82974
rect 333666 47058 333902 47294
rect 333986 47058 334222 47294
rect 333666 46738 333902 46974
rect 333986 46738 334222 46974
rect 333666 11058 333902 11294
rect 333986 11058 334222 11294
rect 333666 10738 333902 10974
rect 333986 10738 334222 10974
rect 341106 708442 341342 708678
rect 341426 708442 341662 708678
rect 341106 708122 341342 708358
rect 341426 708122 341662 708358
rect 341106 666498 341342 666734
rect 341426 666498 341662 666734
rect 341106 666178 341342 666414
rect 341426 666178 341662 666414
rect 341106 630498 341342 630734
rect 341426 630498 341662 630734
rect 341106 630178 341342 630414
rect 341426 630178 341662 630414
rect 341106 594498 341342 594734
rect 341426 594498 341662 594734
rect 341106 594178 341342 594414
rect 341426 594178 341662 594414
rect 341106 558498 341342 558734
rect 341426 558498 341662 558734
rect 341106 558178 341342 558414
rect 341426 558178 341662 558414
rect 341106 522498 341342 522734
rect 341426 522498 341662 522734
rect 341106 522178 341342 522414
rect 341426 522178 341662 522414
rect 341106 486498 341342 486734
rect 341426 486498 341662 486734
rect 341106 486178 341342 486414
rect 341426 486178 341662 486414
rect 341106 450498 341342 450734
rect 341426 450498 341662 450734
rect 341106 450178 341342 450414
rect 341426 450178 341662 450414
rect 341106 414498 341342 414734
rect 341426 414498 341662 414734
rect 341106 414178 341342 414414
rect 341426 414178 341662 414414
rect 341106 378498 341342 378734
rect 341426 378498 341662 378734
rect 341106 378178 341342 378414
rect 341426 378178 341662 378414
rect 341106 342498 341342 342734
rect 341426 342498 341662 342734
rect 341106 342178 341342 342414
rect 341426 342178 341662 342414
rect 341106 306498 341342 306734
rect 341426 306498 341662 306734
rect 341106 306178 341342 306414
rect 341426 306178 341662 306414
rect 341106 270498 341342 270734
rect 341426 270498 341662 270734
rect 341106 270178 341342 270414
rect 341426 270178 341662 270414
rect 341106 234498 341342 234734
rect 341426 234498 341662 234734
rect 341106 234178 341342 234414
rect 341426 234178 341662 234414
rect 341106 198498 341342 198734
rect 341426 198498 341662 198734
rect 341106 198178 341342 198414
rect 341426 198178 341662 198414
rect 341106 162498 341342 162734
rect 341426 162498 341662 162734
rect 341106 162178 341342 162414
rect 341426 162178 341662 162414
rect 341106 126498 341342 126734
rect 341426 126498 341662 126734
rect 341106 126178 341342 126414
rect 341426 126178 341662 126414
rect 337386 86778 337622 87014
rect 337706 86778 337942 87014
rect 337386 86458 337622 86694
rect 337706 86458 337942 86694
rect 337386 50778 337622 51014
rect 337706 50778 337942 51014
rect 337386 50458 337622 50694
rect 337706 50458 337942 50694
rect 337386 14778 337622 15014
rect 337706 14778 337942 15014
rect 337386 14458 337622 14694
rect 337706 14458 337942 14694
rect 333666 -2502 333902 -2266
rect 333986 -2502 334222 -2266
rect 333666 -2822 333902 -2586
rect 333986 -2822 334222 -2586
rect 341106 90498 341342 90734
rect 341426 90498 341662 90734
rect 341106 90178 341342 90414
rect 341426 90178 341662 90414
rect 341106 54498 341342 54734
rect 341426 54498 341662 54734
rect 341106 54178 341342 54414
rect 341426 54178 341662 54414
rect 341106 18498 341342 18734
rect 341426 18498 341662 18734
rect 341106 18178 341342 18414
rect 341426 18178 341662 18414
rect 338902 6342 339138 6578
rect 338350 4302 338586 4538
rect 337386 -3462 337622 -3226
rect 337706 -3462 337942 -3226
rect 337386 -3782 337622 -3546
rect 337706 -3782 337942 -3546
rect 341106 -4422 341342 -4186
rect 341426 -4422 341662 -4186
rect 341106 -4742 341342 -4506
rect 341426 -4742 341662 -4506
rect 344826 709402 345062 709638
rect 345146 709402 345382 709638
rect 344826 709082 345062 709318
rect 345146 709082 345382 709318
rect 344826 670218 345062 670454
rect 345146 670218 345382 670454
rect 344826 669898 345062 670134
rect 345146 669898 345382 670134
rect 344826 634218 345062 634454
rect 345146 634218 345382 634454
rect 344826 633898 345062 634134
rect 345146 633898 345382 634134
rect 344826 598218 345062 598454
rect 345146 598218 345382 598454
rect 344826 597898 345062 598134
rect 345146 597898 345382 598134
rect 344826 562218 345062 562454
rect 345146 562218 345382 562454
rect 344826 561898 345062 562134
rect 345146 561898 345382 562134
rect 344826 526218 345062 526454
rect 345146 526218 345382 526454
rect 344826 525898 345062 526134
rect 345146 525898 345382 526134
rect 344826 490218 345062 490454
rect 345146 490218 345382 490454
rect 344826 489898 345062 490134
rect 345146 489898 345382 490134
rect 344826 454218 345062 454454
rect 345146 454218 345382 454454
rect 344826 453898 345062 454134
rect 345146 453898 345382 454134
rect 344826 418218 345062 418454
rect 345146 418218 345382 418454
rect 344826 417898 345062 418134
rect 345146 417898 345382 418134
rect 344826 382218 345062 382454
rect 345146 382218 345382 382454
rect 344826 381898 345062 382134
rect 345146 381898 345382 382134
rect 344826 346218 345062 346454
rect 345146 346218 345382 346454
rect 344826 345898 345062 346134
rect 345146 345898 345382 346134
rect 344826 310218 345062 310454
rect 345146 310218 345382 310454
rect 344826 309898 345062 310134
rect 345146 309898 345382 310134
rect 344826 274218 345062 274454
rect 345146 274218 345382 274454
rect 344826 273898 345062 274134
rect 345146 273898 345382 274134
rect 344826 238218 345062 238454
rect 345146 238218 345382 238454
rect 344826 237898 345062 238134
rect 345146 237898 345382 238134
rect 344826 202218 345062 202454
rect 345146 202218 345382 202454
rect 344826 201898 345062 202134
rect 345146 201898 345382 202134
rect 344826 166218 345062 166454
rect 345146 166218 345382 166454
rect 344826 165898 345062 166134
rect 345146 165898 345382 166134
rect 344826 130218 345062 130454
rect 345146 130218 345382 130454
rect 344826 129898 345062 130134
rect 345146 129898 345382 130134
rect 344826 94218 345062 94454
rect 345146 94218 345382 94454
rect 344826 93898 345062 94134
rect 345146 93898 345382 94134
rect 344826 58218 345062 58454
rect 345146 58218 345382 58454
rect 344826 57898 345062 58134
rect 345146 57898 345382 58134
rect 344826 22218 345062 22454
rect 345146 22218 345382 22454
rect 344826 21898 345062 22134
rect 345146 21898 345382 22134
rect 344826 -5382 345062 -5146
rect 345146 -5382 345382 -5146
rect 344826 -5702 345062 -5466
rect 345146 -5702 345382 -5466
rect 348546 710362 348782 710598
rect 348866 710362 349102 710598
rect 348546 710042 348782 710278
rect 348866 710042 349102 710278
rect 348546 673938 348782 674174
rect 348866 673938 349102 674174
rect 348546 673618 348782 673854
rect 348866 673618 349102 673854
rect 348546 637938 348782 638174
rect 348866 637938 349102 638174
rect 348546 637618 348782 637854
rect 348866 637618 349102 637854
rect 348546 601938 348782 602174
rect 348866 601938 349102 602174
rect 348546 601618 348782 601854
rect 348866 601618 349102 601854
rect 348546 565938 348782 566174
rect 348866 565938 349102 566174
rect 348546 565618 348782 565854
rect 348866 565618 349102 565854
rect 348546 529938 348782 530174
rect 348866 529938 349102 530174
rect 348546 529618 348782 529854
rect 348866 529618 349102 529854
rect 348546 493938 348782 494174
rect 348866 493938 349102 494174
rect 348546 493618 348782 493854
rect 348866 493618 349102 493854
rect 348546 457938 348782 458174
rect 348866 457938 349102 458174
rect 348546 457618 348782 457854
rect 348866 457618 349102 457854
rect 348546 421938 348782 422174
rect 348866 421938 349102 422174
rect 348546 421618 348782 421854
rect 348866 421618 349102 421854
rect 348546 385938 348782 386174
rect 348866 385938 349102 386174
rect 348546 385618 348782 385854
rect 348866 385618 349102 385854
rect 348546 349938 348782 350174
rect 348866 349938 349102 350174
rect 348546 349618 348782 349854
rect 348866 349618 349102 349854
rect 348546 313938 348782 314174
rect 348866 313938 349102 314174
rect 348546 313618 348782 313854
rect 348866 313618 349102 313854
rect 348546 277938 348782 278174
rect 348866 277938 349102 278174
rect 348546 277618 348782 277854
rect 348866 277618 349102 277854
rect 348546 241938 348782 242174
rect 348866 241938 349102 242174
rect 348546 241618 348782 241854
rect 348866 241618 349102 241854
rect 348546 205938 348782 206174
rect 348866 205938 349102 206174
rect 348546 205618 348782 205854
rect 348866 205618 349102 205854
rect 348546 169938 348782 170174
rect 348866 169938 349102 170174
rect 348546 169618 348782 169854
rect 348866 169618 349102 169854
rect 348546 133938 348782 134174
rect 348866 133938 349102 134174
rect 348546 133618 348782 133854
rect 348866 133618 349102 133854
rect 348546 97938 348782 98174
rect 348866 97938 349102 98174
rect 348546 97618 348782 97854
rect 348866 97618 349102 97854
rect 348546 61938 348782 62174
rect 348866 61938 349102 62174
rect 348546 61618 348782 61854
rect 348866 61618 349102 61854
rect 348546 25938 348782 26174
rect 348866 25938 349102 26174
rect 348546 25618 348782 25854
rect 348866 25618 349102 25854
rect 348546 -6342 348782 -6106
rect 348866 -6342 349102 -6106
rect 348546 -6662 348782 -6426
rect 348866 -6662 349102 -6426
rect 352266 711322 352502 711558
rect 352586 711322 352822 711558
rect 352266 711002 352502 711238
rect 352586 711002 352822 711238
rect 352266 677658 352502 677894
rect 352586 677658 352822 677894
rect 352266 677338 352502 677574
rect 352586 677338 352822 677574
rect 352266 641658 352502 641894
rect 352586 641658 352822 641894
rect 352266 641338 352502 641574
rect 352586 641338 352822 641574
rect 352266 605658 352502 605894
rect 352586 605658 352822 605894
rect 352266 605338 352502 605574
rect 352586 605338 352822 605574
rect 352266 569658 352502 569894
rect 352586 569658 352822 569894
rect 352266 569338 352502 569574
rect 352586 569338 352822 569574
rect 352266 533658 352502 533894
rect 352586 533658 352822 533894
rect 352266 533338 352502 533574
rect 352586 533338 352822 533574
rect 352266 497658 352502 497894
rect 352586 497658 352822 497894
rect 352266 497338 352502 497574
rect 352586 497338 352822 497574
rect 352266 461658 352502 461894
rect 352586 461658 352822 461894
rect 352266 461338 352502 461574
rect 352586 461338 352822 461574
rect 352266 425658 352502 425894
rect 352586 425658 352822 425894
rect 352266 425338 352502 425574
rect 352586 425338 352822 425574
rect 352266 389658 352502 389894
rect 352586 389658 352822 389894
rect 352266 389338 352502 389574
rect 352586 389338 352822 389574
rect 352266 353658 352502 353894
rect 352586 353658 352822 353894
rect 352266 353338 352502 353574
rect 352586 353338 352822 353574
rect 352266 317658 352502 317894
rect 352586 317658 352822 317894
rect 352266 317338 352502 317574
rect 352586 317338 352822 317574
rect 352266 281658 352502 281894
rect 352586 281658 352822 281894
rect 352266 281338 352502 281574
rect 352586 281338 352822 281574
rect 352266 245658 352502 245894
rect 352586 245658 352822 245894
rect 352266 245338 352502 245574
rect 352586 245338 352822 245574
rect 352266 209658 352502 209894
rect 352586 209658 352822 209894
rect 352266 209338 352502 209574
rect 352586 209338 352822 209574
rect 352266 173658 352502 173894
rect 352586 173658 352822 173894
rect 352266 173338 352502 173574
rect 352586 173338 352822 173574
rect 352266 137658 352502 137894
rect 352586 137658 352822 137894
rect 352266 137338 352502 137574
rect 352586 137338 352822 137574
rect 352266 101658 352502 101894
rect 352586 101658 352822 101894
rect 352266 101338 352502 101574
rect 352586 101338 352822 101574
rect 352266 65658 352502 65894
rect 352586 65658 352822 65894
rect 352266 65338 352502 65574
rect 352586 65338 352822 65574
rect 352266 29658 352502 29894
rect 352586 29658 352822 29894
rect 352266 29338 352502 29574
rect 352586 29338 352822 29574
rect 352266 -7302 352502 -7066
rect 352586 -7302 352822 -7066
rect 352266 -7622 352502 -7386
rect 352586 -7622 352822 -7386
rect 362226 704602 362462 704838
rect 362546 704602 362782 704838
rect 362226 704282 362462 704518
rect 362546 704282 362782 704518
rect 362226 687618 362462 687854
rect 362546 687618 362782 687854
rect 362226 687298 362462 687534
rect 362546 687298 362782 687534
rect 362226 651618 362462 651854
rect 362546 651618 362782 651854
rect 362226 651298 362462 651534
rect 362546 651298 362782 651534
rect 362226 615618 362462 615854
rect 362546 615618 362782 615854
rect 362226 615298 362462 615534
rect 362546 615298 362782 615534
rect 362226 579618 362462 579854
rect 362546 579618 362782 579854
rect 362226 579298 362462 579534
rect 362546 579298 362782 579534
rect 362226 543618 362462 543854
rect 362546 543618 362782 543854
rect 362226 543298 362462 543534
rect 362546 543298 362782 543534
rect 362226 507618 362462 507854
rect 362546 507618 362782 507854
rect 362226 507298 362462 507534
rect 362546 507298 362782 507534
rect 362226 471618 362462 471854
rect 362546 471618 362782 471854
rect 362226 471298 362462 471534
rect 362546 471298 362782 471534
rect 362226 435618 362462 435854
rect 362546 435618 362782 435854
rect 362226 435298 362462 435534
rect 362546 435298 362782 435534
rect 362226 399618 362462 399854
rect 362546 399618 362782 399854
rect 362226 399298 362462 399534
rect 362546 399298 362782 399534
rect 362226 363618 362462 363854
rect 362546 363618 362782 363854
rect 362226 363298 362462 363534
rect 362546 363298 362782 363534
rect 362226 327618 362462 327854
rect 362546 327618 362782 327854
rect 362226 327298 362462 327534
rect 362546 327298 362782 327534
rect 362226 291618 362462 291854
rect 362546 291618 362782 291854
rect 362226 291298 362462 291534
rect 362546 291298 362782 291534
rect 362226 255618 362462 255854
rect 362546 255618 362782 255854
rect 362226 255298 362462 255534
rect 362546 255298 362782 255534
rect 362226 219618 362462 219854
rect 362546 219618 362782 219854
rect 362226 219298 362462 219534
rect 362546 219298 362782 219534
rect 362226 183618 362462 183854
rect 362546 183618 362782 183854
rect 362226 183298 362462 183534
rect 362546 183298 362782 183534
rect 362226 147618 362462 147854
rect 362546 147618 362782 147854
rect 362226 147298 362462 147534
rect 362546 147298 362782 147534
rect 362226 111618 362462 111854
rect 362546 111618 362782 111854
rect 362226 111298 362462 111534
rect 362546 111298 362782 111534
rect 362226 75618 362462 75854
rect 362546 75618 362782 75854
rect 362226 75298 362462 75534
rect 362546 75298 362782 75534
rect 362226 39618 362462 39854
rect 362546 39618 362782 39854
rect 362226 39298 362462 39534
rect 362546 39298 362782 39534
rect 362226 3618 362462 3854
rect 362546 3618 362782 3854
rect 362226 3298 362462 3534
rect 362546 3298 362782 3534
rect 362226 -582 362462 -346
rect 362546 -582 362782 -346
rect 362226 -902 362462 -666
rect 362546 -902 362782 -666
rect 365946 705562 366182 705798
rect 366266 705562 366502 705798
rect 365946 705242 366182 705478
rect 366266 705242 366502 705478
rect 365946 691338 366182 691574
rect 366266 691338 366502 691574
rect 365946 691018 366182 691254
rect 366266 691018 366502 691254
rect 365946 655338 366182 655574
rect 366266 655338 366502 655574
rect 365946 655018 366182 655254
rect 366266 655018 366502 655254
rect 365946 619338 366182 619574
rect 366266 619338 366502 619574
rect 365946 619018 366182 619254
rect 366266 619018 366502 619254
rect 365946 583338 366182 583574
rect 366266 583338 366502 583574
rect 365946 583018 366182 583254
rect 366266 583018 366502 583254
rect 365946 547338 366182 547574
rect 366266 547338 366502 547574
rect 365946 547018 366182 547254
rect 366266 547018 366502 547254
rect 365946 511338 366182 511574
rect 366266 511338 366502 511574
rect 365946 511018 366182 511254
rect 366266 511018 366502 511254
rect 365946 475338 366182 475574
rect 366266 475338 366502 475574
rect 365946 475018 366182 475254
rect 366266 475018 366502 475254
rect 365946 439338 366182 439574
rect 366266 439338 366502 439574
rect 365946 439018 366182 439254
rect 366266 439018 366502 439254
rect 365946 403338 366182 403574
rect 366266 403338 366502 403574
rect 365946 403018 366182 403254
rect 366266 403018 366502 403254
rect 365946 367338 366182 367574
rect 366266 367338 366502 367574
rect 365946 367018 366182 367254
rect 366266 367018 366502 367254
rect 365946 331338 366182 331574
rect 366266 331338 366502 331574
rect 365946 331018 366182 331254
rect 366266 331018 366502 331254
rect 365946 295338 366182 295574
rect 366266 295338 366502 295574
rect 365946 295018 366182 295254
rect 366266 295018 366502 295254
rect 365946 259338 366182 259574
rect 366266 259338 366502 259574
rect 365946 259018 366182 259254
rect 366266 259018 366502 259254
rect 365946 223338 366182 223574
rect 366266 223338 366502 223574
rect 365946 223018 366182 223254
rect 366266 223018 366502 223254
rect 365946 187338 366182 187574
rect 366266 187338 366502 187574
rect 365946 187018 366182 187254
rect 366266 187018 366502 187254
rect 365946 151338 366182 151574
rect 366266 151338 366502 151574
rect 365946 151018 366182 151254
rect 366266 151018 366502 151254
rect 365946 115338 366182 115574
rect 366266 115338 366502 115574
rect 365946 115018 366182 115254
rect 366266 115018 366502 115254
rect 365946 79338 366182 79574
rect 366266 79338 366502 79574
rect 365946 79018 366182 79254
rect 366266 79018 366502 79254
rect 365946 43338 366182 43574
rect 366266 43338 366502 43574
rect 365946 43018 366182 43254
rect 366266 43018 366502 43254
rect 365946 7338 366182 7574
rect 366266 7338 366502 7574
rect 365946 7018 366182 7254
rect 366266 7018 366502 7254
rect 365946 -1542 366182 -1306
rect 366266 -1542 366502 -1306
rect 365946 -1862 366182 -1626
rect 366266 -1862 366502 -1626
rect 369666 706522 369902 706758
rect 369986 706522 370222 706758
rect 369666 706202 369902 706438
rect 369986 706202 370222 706438
rect 369666 695058 369902 695294
rect 369986 695058 370222 695294
rect 369666 694738 369902 694974
rect 369986 694738 370222 694974
rect 369666 659058 369902 659294
rect 369986 659058 370222 659294
rect 369666 658738 369902 658974
rect 369986 658738 370222 658974
rect 369666 623058 369902 623294
rect 369986 623058 370222 623294
rect 369666 622738 369902 622974
rect 369986 622738 370222 622974
rect 369666 587058 369902 587294
rect 369986 587058 370222 587294
rect 369666 586738 369902 586974
rect 369986 586738 370222 586974
rect 369666 551058 369902 551294
rect 369986 551058 370222 551294
rect 369666 550738 369902 550974
rect 369986 550738 370222 550974
rect 369666 515058 369902 515294
rect 369986 515058 370222 515294
rect 369666 514738 369902 514974
rect 369986 514738 370222 514974
rect 369666 479058 369902 479294
rect 369986 479058 370222 479294
rect 369666 478738 369902 478974
rect 369986 478738 370222 478974
rect 369666 443058 369902 443294
rect 369986 443058 370222 443294
rect 369666 442738 369902 442974
rect 369986 442738 370222 442974
rect 369666 407058 369902 407294
rect 369986 407058 370222 407294
rect 369666 406738 369902 406974
rect 369986 406738 370222 406974
rect 369666 371058 369902 371294
rect 369986 371058 370222 371294
rect 369666 370738 369902 370974
rect 369986 370738 370222 370974
rect 369666 335058 369902 335294
rect 369986 335058 370222 335294
rect 369666 334738 369902 334974
rect 369986 334738 370222 334974
rect 369666 299058 369902 299294
rect 369986 299058 370222 299294
rect 369666 298738 369902 298974
rect 369986 298738 370222 298974
rect 369666 263058 369902 263294
rect 369986 263058 370222 263294
rect 369666 262738 369902 262974
rect 369986 262738 370222 262974
rect 369666 227058 369902 227294
rect 369986 227058 370222 227294
rect 369666 226738 369902 226974
rect 369986 226738 370222 226974
rect 369666 191058 369902 191294
rect 369986 191058 370222 191294
rect 369666 190738 369902 190974
rect 369986 190738 370222 190974
rect 369666 155058 369902 155294
rect 369986 155058 370222 155294
rect 369666 154738 369902 154974
rect 369986 154738 370222 154974
rect 369666 119058 369902 119294
rect 369986 119058 370222 119294
rect 369666 118738 369902 118974
rect 369986 118738 370222 118974
rect 369666 83058 369902 83294
rect 369986 83058 370222 83294
rect 369666 82738 369902 82974
rect 369986 82738 370222 82974
rect 369666 47058 369902 47294
rect 369986 47058 370222 47294
rect 369666 46738 369902 46974
rect 369986 46738 370222 46974
rect 369666 11058 369902 11294
rect 369986 11058 370222 11294
rect 369666 10738 369902 10974
rect 369986 10738 370222 10974
rect 369666 -2502 369902 -2266
rect 369986 -2502 370222 -2266
rect 369666 -2822 369902 -2586
rect 369986 -2822 370222 -2586
rect 373386 707482 373622 707718
rect 373706 707482 373942 707718
rect 373386 707162 373622 707398
rect 373706 707162 373942 707398
rect 373386 698778 373622 699014
rect 373706 698778 373942 699014
rect 373386 698458 373622 698694
rect 373706 698458 373942 698694
rect 373386 662778 373622 663014
rect 373706 662778 373942 663014
rect 373386 662458 373622 662694
rect 373706 662458 373942 662694
rect 373386 626778 373622 627014
rect 373706 626778 373942 627014
rect 373386 626458 373622 626694
rect 373706 626458 373942 626694
rect 373386 590778 373622 591014
rect 373706 590778 373942 591014
rect 373386 590458 373622 590694
rect 373706 590458 373942 590694
rect 373386 554778 373622 555014
rect 373706 554778 373942 555014
rect 373386 554458 373622 554694
rect 373706 554458 373942 554694
rect 373386 518778 373622 519014
rect 373706 518778 373942 519014
rect 373386 518458 373622 518694
rect 373706 518458 373942 518694
rect 373386 482778 373622 483014
rect 373706 482778 373942 483014
rect 373386 482458 373622 482694
rect 373706 482458 373942 482694
rect 373386 446778 373622 447014
rect 373706 446778 373942 447014
rect 373386 446458 373622 446694
rect 373706 446458 373942 446694
rect 373386 410778 373622 411014
rect 373706 410778 373942 411014
rect 373386 410458 373622 410694
rect 373706 410458 373942 410694
rect 373386 374778 373622 375014
rect 373706 374778 373942 375014
rect 373386 374458 373622 374694
rect 373706 374458 373942 374694
rect 373386 338778 373622 339014
rect 373706 338778 373942 339014
rect 373386 338458 373622 338694
rect 373706 338458 373942 338694
rect 373386 302778 373622 303014
rect 373706 302778 373942 303014
rect 373386 302458 373622 302694
rect 373706 302458 373942 302694
rect 373386 266778 373622 267014
rect 373706 266778 373942 267014
rect 373386 266458 373622 266694
rect 373706 266458 373942 266694
rect 373386 230778 373622 231014
rect 373706 230778 373942 231014
rect 373386 230458 373622 230694
rect 373706 230458 373942 230694
rect 373386 194778 373622 195014
rect 373706 194778 373942 195014
rect 373386 194458 373622 194694
rect 373706 194458 373942 194694
rect 373386 158778 373622 159014
rect 373706 158778 373942 159014
rect 373386 158458 373622 158694
rect 373706 158458 373942 158694
rect 373386 122778 373622 123014
rect 373706 122778 373942 123014
rect 373386 122458 373622 122694
rect 373706 122458 373942 122694
rect 373386 86778 373622 87014
rect 373706 86778 373942 87014
rect 373386 86458 373622 86694
rect 373706 86458 373942 86694
rect 373386 50778 373622 51014
rect 373706 50778 373942 51014
rect 373386 50458 373622 50694
rect 373706 50458 373942 50694
rect 373386 14778 373622 15014
rect 373706 14778 373942 15014
rect 373386 14458 373622 14694
rect 373706 14458 373942 14694
rect 373386 -3462 373622 -3226
rect 373706 -3462 373942 -3226
rect 373386 -3782 373622 -3546
rect 373706 -3782 373942 -3546
rect 377106 708442 377342 708678
rect 377426 708442 377662 708678
rect 377106 708122 377342 708358
rect 377426 708122 377662 708358
rect 377106 666498 377342 666734
rect 377426 666498 377662 666734
rect 377106 666178 377342 666414
rect 377426 666178 377662 666414
rect 377106 630498 377342 630734
rect 377426 630498 377662 630734
rect 377106 630178 377342 630414
rect 377426 630178 377662 630414
rect 377106 594498 377342 594734
rect 377426 594498 377662 594734
rect 377106 594178 377342 594414
rect 377426 594178 377662 594414
rect 377106 558498 377342 558734
rect 377426 558498 377662 558734
rect 377106 558178 377342 558414
rect 377426 558178 377662 558414
rect 377106 522498 377342 522734
rect 377426 522498 377662 522734
rect 377106 522178 377342 522414
rect 377426 522178 377662 522414
rect 377106 486498 377342 486734
rect 377426 486498 377662 486734
rect 377106 486178 377342 486414
rect 377426 486178 377662 486414
rect 377106 450498 377342 450734
rect 377426 450498 377662 450734
rect 377106 450178 377342 450414
rect 377426 450178 377662 450414
rect 377106 414498 377342 414734
rect 377426 414498 377662 414734
rect 377106 414178 377342 414414
rect 377426 414178 377662 414414
rect 377106 378498 377342 378734
rect 377426 378498 377662 378734
rect 377106 378178 377342 378414
rect 377426 378178 377662 378414
rect 377106 342498 377342 342734
rect 377426 342498 377662 342734
rect 377106 342178 377342 342414
rect 377426 342178 377662 342414
rect 377106 306498 377342 306734
rect 377426 306498 377662 306734
rect 377106 306178 377342 306414
rect 377426 306178 377662 306414
rect 377106 270498 377342 270734
rect 377426 270498 377662 270734
rect 377106 270178 377342 270414
rect 377426 270178 377662 270414
rect 377106 234498 377342 234734
rect 377426 234498 377662 234734
rect 377106 234178 377342 234414
rect 377426 234178 377662 234414
rect 377106 198498 377342 198734
rect 377426 198498 377662 198734
rect 377106 198178 377342 198414
rect 377426 198178 377662 198414
rect 377106 162498 377342 162734
rect 377426 162498 377662 162734
rect 377106 162178 377342 162414
rect 377426 162178 377662 162414
rect 377106 126498 377342 126734
rect 377426 126498 377662 126734
rect 377106 126178 377342 126414
rect 377426 126178 377662 126414
rect 377106 90498 377342 90734
rect 377426 90498 377662 90734
rect 377106 90178 377342 90414
rect 377426 90178 377662 90414
rect 377106 54498 377342 54734
rect 377426 54498 377662 54734
rect 377106 54178 377342 54414
rect 377426 54178 377662 54414
rect 377106 18498 377342 18734
rect 377426 18498 377662 18734
rect 377106 18178 377342 18414
rect 377426 18178 377662 18414
rect 377106 -4422 377342 -4186
rect 377426 -4422 377662 -4186
rect 377106 -4742 377342 -4506
rect 377426 -4742 377662 -4506
rect 380826 709402 381062 709638
rect 381146 709402 381382 709638
rect 380826 709082 381062 709318
rect 381146 709082 381382 709318
rect 380826 670218 381062 670454
rect 381146 670218 381382 670454
rect 380826 669898 381062 670134
rect 381146 669898 381382 670134
rect 380826 634218 381062 634454
rect 381146 634218 381382 634454
rect 380826 633898 381062 634134
rect 381146 633898 381382 634134
rect 380826 598218 381062 598454
rect 381146 598218 381382 598454
rect 380826 597898 381062 598134
rect 381146 597898 381382 598134
rect 380826 562218 381062 562454
rect 381146 562218 381382 562454
rect 380826 561898 381062 562134
rect 381146 561898 381382 562134
rect 380826 526218 381062 526454
rect 381146 526218 381382 526454
rect 380826 525898 381062 526134
rect 381146 525898 381382 526134
rect 380826 490218 381062 490454
rect 381146 490218 381382 490454
rect 380826 489898 381062 490134
rect 381146 489898 381382 490134
rect 380826 454218 381062 454454
rect 381146 454218 381382 454454
rect 380826 453898 381062 454134
rect 381146 453898 381382 454134
rect 380826 418218 381062 418454
rect 381146 418218 381382 418454
rect 380826 417898 381062 418134
rect 381146 417898 381382 418134
rect 380826 382218 381062 382454
rect 381146 382218 381382 382454
rect 380826 381898 381062 382134
rect 381146 381898 381382 382134
rect 380826 346218 381062 346454
rect 381146 346218 381382 346454
rect 380826 345898 381062 346134
rect 381146 345898 381382 346134
rect 380826 310218 381062 310454
rect 381146 310218 381382 310454
rect 380826 309898 381062 310134
rect 381146 309898 381382 310134
rect 380826 274218 381062 274454
rect 381146 274218 381382 274454
rect 380826 273898 381062 274134
rect 381146 273898 381382 274134
rect 380826 238218 381062 238454
rect 381146 238218 381382 238454
rect 380826 237898 381062 238134
rect 381146 237898 381382 238134
rect 380826 202218 381062 202454
rect 381146 202218 381382 202454
rect 380826 201898 381062 202134
rect 381146 201898 381382 202134
rect 380826 166218 381062 166454
rect 381146 166218 381382 166454
rect 380826 165898 381062 166134
rect 381146 165898 381382 166134
rect 380826 130218 381062 130454
rect 381146 130218 381382 130454
rect 380826 129898 381062 130134
rect 381146 129898 381382 130134
rect 380826 94218 381062 94454
rect 381146 94218 381382 94454
rect 380826 93898 381062 94134
rect 381146 93898 381382 94134
rect 380826 58218 381062 58454
rect 381146 58218 381382 58454
rect 380826 57898 381062 58134
rect 381146 57898 381382 58134
rect 380826 22218 381062 22454
rect 381146 22218 381382 22454
rect 380826 21898 381062 22134
rect 381146 21898 381382 22134
rect 380826 -5382 381062 -5146
rect 381146 -5382 381382 -5146
rect 380826 -5702 381062 -5466
rect 381146 -5702 381382 -5466
rect 384546 710362 384782 710598
rect 384866 710362 385102 710598
rect 384546 710042 384782 710278
rect 384866 710042 385102 710278
rect 384546 673938 384782 674174
rect 384866 673938 385102 674174
rect 384546 673618 384782 673854
rect 384866 673618 385102 673854
rect 384546 637938 384782 638174
rect 384866 637938 385102 638174
rect 384546 637618 384782 637854
rect 384866 637618 385102 637854
rect 384546 601938 384782 602174
rect 384866 601938 385102 602174
rect 384546 601618 384782 601854
rect 384866 601618 385102 601854
rect 384546 565938 384782 566174
rect 384866 565938 385102 566174
rect 384546 565618 384782 565854
rect 384866 565618 385102 565854
rect 384546 529938 384782 530174
rect 384866 529938 385102 530174
rect 384546 529618 384782 529854
rect 384866 529618 385102 529854
rect 384546 493938 384782 494174
rect 384866 493938 385102 494174
rect 384546 493618 384782 493854
rect 384866 493618 385102 493854
rect 384546 457938 384782 458174
rect 384866 457938 385102 458174
rect 384546 457618 384782 457854
rect 384866 457618 385102 457854
rect 384546 421938 384782 422174
rect 384866 421938 385102 422174
rect 384546 421618 384782 421854
rect 384866 421618 385102 421854
rect 384546 385938 384782 386174
rect 384866 385938 385102 386174
rect 384546 385618 384782 385854
rect 384866 385618 385102 385854
rect 384546 349938 384782 350174
rect 384866 349938 385102 350174
rect 384546 349618 384782 349854
rect 384866 349618 385102 349854
rect 384546 313938 384782 314174
rect 384866 313938 385102 314174
rect 384546 313618 384782 313854
rect 384866 313618 385102 313854
rect 384546 277938 384782 278174
rect 384866 277938 385102 278174
rect 384546 277618 384782 277854
rect 384866 277618 385102 277854
rect 384546 241938 384782 242174
rect 384866 241938 385102 242174
rect 384546 241618 384782 241854
rect 384866 241618 385102 241854
rect 384546 205938 384782 206174
rect 384866 205938 385102 206174
rect 384546 205618 384782 205854
rect 384866 205618 385102 205854
rect 384546 169938 384782 170174
rect 384866 169938 385102 170174
rect 384546 169618 384782 169854
rect 384866 169618 385102 169854
rect 384546 133938 384782 134174
rect 384866 133938 385102 134174
rect 384546 133618 384782 133854
rect 384866 133618 385102 133854
rect 384546 97938 384782 98174
rect 384866 97938 385102 98174
rect 384546 97618 384782 97854
rect 384866 97618 385102 97854
rect 384546 61938 384782 62174
rect 384866 61938 385102 62174
rect 384546 61618 384782 61854
rect 384866 61618 385102 61854
rect 384546 25938 384782 26174
rect 384866 25938 385102 26174
rect 384546 25618 384782 25854
rect 384866 25618 385102 25854
rect 384546 -6342 384782 -6106
rect 384866 -6342 385102 -6106
rect 384546 -6662 384782 -6426
rect 384866 -6662 385102 -6426
rect 388266 711322 388502 711558
rect 388586 711322 388822 711558
rect 388266 711002 388502 711238
rect 388586 711002 388822 711238
rect 388266 677658 388502 677894
rect 388586 677658 388822 677894
rect 388266 677338 388502 677574
rect 388586 677338 388822 677574
rect 388266 641658 388502 641894
rect 388586 641658 388822 641894
rect 388266 641338 388502 641574
rect 388586 641338 388822 641574
rect 388266 605658 388502 605894
rect 388586 605658 388822 605894
rect 388266 605338 388502 605574
rect 388586 605338 388822 605574
rect 388266 569658 388502 569894
rect 388586 569658 388822 569894
rect 388266 569338 388502 569574
rect 388586 569338 388822 569574
rect 388266 533658 388502 533894
rect 388586 533658 388822 533894
rect 388266 533338 388502 533574
rect 388586 533338 388822 533574
rect 388266 497658 388502 497894
rect 388586 497658 388822 497894
rect 388266 497338 388502 497574
rect 388586 497338 388822 497574
rect 388266 461658 388502 461894
rect 388586 461658 388822 461894
rect 388266 461338 388502 461574
rect 388586 461338 388822 461574
rect 388266 425658 388502 425894
rect 388586 425658 388822 425894
rect 388266 425338 388502 425574
rect 388586 425338 388822 425574
rect 388266 389658 388502 389894
rect 388586 389658 388822 389894
rect 388266 389338 388502 389574
rect 388586 389338 388822 389574
rect 388266 353658 388502 353894
rect 388586 353658 388822 353894
rect 388266 353338 388502 353574
rect 388586 353338 388822 353574
rect 388266 317658 388502 317894
rect 388586 317658 388822 317894
rect 388266 317338 388502 317574
rect 388586 317338 388822 317574
rect 388266 281658 388502 281894
rect 388586 281658 388822 281894
rect 388266 281338 388502 281574
rect 388586 281338 388822 281574
rect 388266 245658 388502 245894
rect 388586 245658 388822 245894
rect 388266 245338 388502 245574
rect 388586 245338 388822 245574
rect 388266 209658 388502 209894
rect 388586 209658 388822 209894
rect 388266 209338 388502 209574
rect 388586 209338 388822 209574
rect 388266 173658 388502 173894
rect 388586 173658 388822 173894
rect 388266 173338 388502 173574
rect 388586 173338 388822 173574
rect 388266 137658 388502 137894
rect 388586 137658 388822 137894
rect 388266 137338 388502 137574
rect 388586 137338 388822 137574
rect 388266 101658 388502 101894
rect 388586 101658 388822 101894
rect 388266 101338 388502 101574
rect 388586 101338 388822 101574
rect 388266 65658 388502 65894
rect 388586 65658 388822 65894
rect 388266 65338 388502 65574
rect 388586 65338 388822 65574
rect 388266 29658 388502 29894
rect 388586 29658 388822 29894
rect 388266 29338 388502 29574
rect 388586 29338 388822 29574
rect 388266 -7302 388502 -7066
rect 388586 -7302 388822 -7066
rect 388266 -7622 388502 -7386
rect 388586 -7622 388822 -7386
rect 398226 704602 398462 704838
rect 398546 704602 398782 704838
rect 398226 704282 398462 704518
rect 398546 704282 398782 704518
rect 398226 687618 398462 687854
rect 398546 687618 398782 687854
rect 398226 687298 398462 687534
rect 398546 687298 398782 687534
rect 398226 651618 398462 651854
rect 398546 651618 398782 651854
rect 398226 651298 398462 651534
rect 398546 651298 398782 651534
rect 398226 615618 398462 615854
rect 398546 615618 398782 615854
rect 398226 615298 398462 615534
rect 398546 615298 398782 615534
rect 398226 579618 398462 579854
rect 398546 579618 398782 579854
rect 398226 579298 398462 579534
rect 398546 579298 398782 579534
rect 398226 543618 398462 543854
rect 398546 543618 398782 543854
rect 398226 543298 398462 543534
rect 398546 543298 398782 543534
rect 398226 507618 398462 507854
rect 398546 507618 398782 507854
rect 398226 507298 398462 507534
rect 398546 507298 398782 507534
rect 398226 471618 398462 471854
rect 398546 471618 398782 471854
rect 398226 471298 398462 471534
rect 398546 471298 398782 471534
rect 398226 435618 398462 435854
rect 398546 435618 398782 435854
rect 398226 435298 398462 435534
rect 398546 435298 398782 435534
rect 398226 399618 398462 399854
rect 398546 399618 398782 399854
rect 398226 399298 398462 399534
rect 398546 399298 398782 399534
rect 398226 363618 398462 363854
rect 398546 363618 398782 363854
rect 398226 363298 398462 363534
rect 398546 363298 398782 363534
rect 398226 327618 398462 327854
rect 398546 327618 398782 327854
rect 398226 327298 398462 327534
rect 398546 327298 398782 327534
rect 398226 291618 398462 291854
rect 398546 291618 398782 291854
rect 398226 291298 398462 291534
rect 398546 291298 398782 291534
rect 398226 255618 398462 255854
rect 398546 255618 398782 255854
rect 398226 255298 398462 255534
rect 398546 255298 398782 255534
rect 398226 219618 398462 219854
rect 398546 219618 398782 219854
rect 398226 219298 398462 219534
rect 398546 219298 398782 219534
rect 398226 183618 398462 183854
rect 398546 183618 398782 183854
rect 398226 183298 398462 183534
rect 398546 183298 398782 183534
rect 398226 147618 398462 147854
rect 398546 147618 398782 147854
rect 398226 147298 398462 147534
rect 398546 147298 398782 147534
rect 398226 111618 398462 111854
rect 398546 111618 398782 111854
rect 398226 111298 398462 111534
rect 398546 111298 398782 111534
rect 398226 75618 398462 75854
rect 398546 75618 398782 75854
rect 398226 75298 398462 75534
rect 398546 75298 398782 75534
rect 398226 39618 398462 39854
rect 398546 39618 398782 39854
rect 398226 39298 398462 39534
rect 398546 39298 398782 39534
rect 398226 3618 398462 3854
rect 398546 3618 398782 3854
rect 398226 3298 398462 3534
rect 398546 3298 398782 3534
rect 398226 -582 398462 -346
rect 398546 -582 398782 -346
rect 398226 -902 398462 -666
rect 398546 -902 398782 -666
rect 401946 705562 402182 705798
rect 402266 705562 402502 705798
rect 401946 705242 402182 705478
rect 402266 705242 402502 705478
rect 401946 691338 402182 691574
rect 402266 691338 402502 691574
rect 401946 691018 402182 691254
rect 402266 691018 402502 691254
rect 401946 655338 402182 655574
rect 402266 655338 402502 655574
rect 401946 655018 402182 655254
rect 402266 655018 402502 655254
rect 401946 619338 402182 619574
rect 402266 619338 402502 619574
rect 401946 619018 402182 619254
rect 402266 619018 402502 619254
rect 401946 583338 402182 583574
rect 402266 583338 402502 583574
rect 401946 583018 402182 583254
rect 402266 583018 402502 583254
rect 401946 547338 402182 547574
rect 402266 547338 402502 547574
rect 401946 547018 402182 547254
rect 402266 547018 402502 547254
rect 401946 511338 402182 511574
rect 402266 511338 402502 511574
rect 401946 511018 402182 511254
rect 402266 511018 402502 511254
rect 401946 475338 402182 475574
rect 402266 475338 402502 475574
rect 401946 475018 402182 475254
rect 402266 475018 402502 475254
rect 401946 439338 402182 439574
rect 402266 439338 402502 439574
rect 401946 439018 402182 439254
rect 402266 439018 402502 439254
rect 401946 403338 402182 403574
rect 402266 403338 402502 403574
rect 401946 403018 402182 403254
rect 402266 403018 402502 403254
rect 401946 367338 402182 367574
rect 402266 367338 402502 367574
rect 401946 367018 402182 367254
rect 402266 367018 402502 367254
rect 401946 331338 402182 331574
rect 402266 331338 402502 331574
rect 401946 331018 402182 331254
rect 402266 331018 402502 331254
rect 401946 295338 402182 295574
rect 402266 295338 402502 295574
rect 401946 295018 402182 295254
rect 402266 295018 402502 295254
rect 401946 259338 402182 259574
rect 402266 259338 402502 259574
rect 401946 259018 402182 259254
rect 402266 259018 402502 259254
rect 401946 223338 402182 223574
rect 402266 223338 402502 223574
rect 401946 223018 402182 223254
rect 402266 223018 402502 223254
rect 401946 187338 402182 187574
rect 402266 187338 402502 187574
rect 401946 187018 402182 187254
rect 402266 187018 402502 187254
rect 401946 151338 402182 151574
rect 402266 151338 402502 151574
rect 401946 151018 402182 151254
rect 402266 151018 402502 151254
rect 401946 115338 402182 115574
rect 402266 115338 402502 115574
rect 401946 115018 402182 115254
rect 402266 115018 402502 115254
rect 405666 706522 405902 706758
rect 405986 706522 406222 706758
rect 405666 706202 405902 706438
rect 405986 706202 406222 706438
rect 405666 695058 405902 695294
rect 405986 695058 406222 695294
rect 405666 694738 405902 694974
rect 405986 694738 406222 694974
rect 405666 659058 405902 659294
rect 405986 659058 406222 659294
rect 405666 658738 405902 658974
rect 405986 658738 406222 658974
rect 405666 623058 405902 623294
rect 405986 623058 406222 623294
rect 405666 622738 405902 622974
rect 405986 622738 406222 622974
rect 405666 587058 405902 587294
rect 405986 587058 406222 587294
rect 405666 586738 405902 586974
rect 405986 586738 406222 586974
rect 405666 551058 405902 551294
rect 405986 551058 406222 551294
rect 405666 550738 405902 550974
rect 405986 550738 406222 550974
rect 405666 515058 405902 515294
rect 405986 515058 406222 515294
rect 405666 514738 405902 514974
rect 405986 514738 406222 514974
rect 405666 479058 405902 479294
rect 405986 479058 406222 479294
rect 405666 478738 405902 478974
rect 405986 478738 406222 478974
rect 405666 443058 405902 443294
rect 405986 443058 406222 443294
rect 405666 442738 405902 442974
rect 405986 442738 406222 442974
rect 405666 407058 405902 407294
rect 405986 407058 406222 407294
rect 405666 406738 405902 406974
rect 405986 406738 406222 406974
rect 405666 371058 405902 371294
rect 405986 371058 406222 371294
rect 405666 370738 405902 370974
rect 405986 370738 406222 370974
rect 405666 335058 405902 335294
rect 405986 335058 406222 335294
rect 405666 334738 405902 334974
rect 405986 334738 406222 334974
rect 405666 299058 405902 299294
rect 405986 299058 406222 299294
rect 405666 298738 405902 298974
rect 405986 298738 406222 298974
rect 405666 263058 405902 263294
rect 405986 263058 406222 263294
rect 405666 262738 405902 262974
rect 405986 262738 406222 262974
rect 405666 227058 405902 227294
rect 405986 227058 406222 227294
rect 405666 226738 405902 226974
rect 405986 226738 406222 226974
rect 405666 191058 405902 191294
rect 405986 191058 406222 191294
rect 405666 190738 405902 190974
rect 405986 190738 406222 190974
rect 405666 155058 405902 155294
rect 405986 155058 406222 155294
rect 405666 154738 405902 154974
rect 405986 154738 406222 154974
rect 405666 119058 405902 119294
rect 405986 119058 406222 119294
rect 405666 118738 405902 118974
rect 405986 118738 406222 118974
rect 404250 111618 404486 111854
rect 404250 111298 404486 111534
rect 401946 79338 402182 79574
rect 402266 79338 402502 79574
rect 401946 79018 402182 79254
rect 402266 79018 402502 79254
rect 401946 43338 402182 43574
rect 402266 43338 402502 43574
rect 401946 43018 402182 43254
rect 402266 43018 402502 43254
rect 401946 7338 402182 7574
rect 402266 7338 402502 7574
rect 401946 7018 402182 7254
rect 402266 7018 402502 7254
rect 401946 -1542 402182 -1306
rect 402266 -1542 402502 -1306
rect 401946 -1862 402182 -1626
rect 402266 -1862 402502 -1626
rect 405666 83058 405902 83294
rect 405986 83058 406222 83294
rect 405666 82738 405902 82974
rect 405986 82738 406222 82974
rect 409386 707482 409622 707718
rect 409706 707482 409942 707718
rect 409386 707162 409622 707398
rect 409706 707162 409942 707398
rect 409386 698778 409622 699014
rect 409706 698778 409942 699014
rect 409386 698458 409622 698694
rect 409706 698458 409942 698694
rect 409386 662778 409622 663014
rect 409706 662778 409942 663014
rect 409386 662458 409622 662694
rect 409706 662458 409942 662694
rect 409386 626778 409622 627014
rect 409706 626778 409942 627014
rect 409386 626458 409622 626694
rect 409706 626458 409942 626694
rect 409386 590778 409622 591014
rect 409706 590778 409942 591014
rect 409386 590458 409622 590694
rect 409706 590458 409942 590694
rect 409386 554778 409622 555014
rect 409706 554778 409942 555014
rect 409386 554458 409622 554694
rect 409706 554458 409942 554694
rect 409386 518778 409622 519014
rect 409706 518778 409942 519014
rect 409386 518458 409622 518694
rect 409706 518458 409942 518694
rect 409386 482778 409622 483014
rect 409706 482778 409942 483014
rect 409386 482458 409622 482694
rect 409706 482458 409942 482694
rect 409386 446778 409622 447014
rect 409706 446778 409942 447014
rect 409386 446458 409622 446694
rect 409706 446458 409942 446694
rect 409386 410778 409622 411014
rect 409706 410778 409942 411014
rect 409386 410458 409622 410694
rect 409706 410458 409942 410694
rect 409386 374778 409622 375014
rect 409706 374778 409942 375014
rect 409386 374458 409622 374694
rect 409706 374458 409942 374694
rect 409386 338778 409622 339014
rect 409706 338778 409942 339014
rect 409386 338458 409622 338694
rect 409706 338458 409942 338694
rect 409386 302778 409622 303014
rect 409706 302778 409942 303014
rect 409386 302458 409622 302694
rect 409706 302458 409942 302694
rect 409386 266778 409622 267014
rect 409706 266778 409942 267014
rect 409386 266458 409622 266694
rect 409706 266458 409942 266694
rect 409386 230778 409622 231014
rect 409706 230778 409942 231014
rect 409386 230458 409622 230694
rect 409706 230458 409942 230694
rect 409386 194778 409622 195014
rect 409706 194778 409942 195014
rect 409386 194458 409622 194694
rect 409706 194458 409942 194694
rect 409386 158778 409622 159014
rect 409706 158778 409942 159014
rect 409386 158458 409622 158694
rect 409706 158458 409942 158694
rect 413106 708442 413342 708678
rect 413426 708442 413662 708678
rect 413106 708122 413342 708358
rect 413426 708122 413662 708358
rect 413106 666498 413342 666734
rect 413426 666498 413662 666734
rect 413106 666178 413342 666414
rect 413426 666178 413662 666414
rect 413106 630498 413342 630734
rect 413426 630498 413662 630734
rect 413106 630178 413342 630414
rect 413426 630178 413662 630414
rect 413106 594498 413342 594734
rect 413426 594498 413662 594734
rect 413106 594178 413342 594414
rect 413426 594178 413662 594414
rect 413106 558498 413342 558734
rect 413426 558498 413662 558734
rect 413106 558178 413342 558414
rect 413426 558178 413662 558414
rect 413106 522498 413342 522734
rect 413426 522498 413662 522734
rect 413106 522178 413342 522414
rect 413426 522178 413662 522414
rect 413106 486498 413342 486734
rect 413426 486498 413662 486734
rect 413106 486178 413342 486414
rect 413426 486178 413662 486414
rect 413106 450498 413342 450734
rect 413426 450498 413662 450734
rect 413106 450178 413342 450414
rect 413426 450178 413662 450414
rect 413106 414498 413342 414734
rect 413426 414498 413662 414734
rect 413106 414178 413342 414414
rect 413426 414178 413662 414414
rect 413106 378498 413342 378734
rect 413426 378498 413662 378734
rect 413106 378178 413342 378414
rect 413426 378178 413662 378414
rect 413106 342498 413342 342734
rect 413426 342498 413662 342734
rect 413106 342178 413342 342414
rect 413426 342178 413662 342414
rect 413106 306498 413342 306734
rect 413426 306498 413662 306734
rect 413106 306178 413342 306414
rect 413426 306178 413662 306414
rect 413106 270498 413342 270734
rect 413426 270498 413662 270734
rect 413106 270178 413342 270414
rect 413426 270178 413662 270414
rect 413106 234498 413342 234734
rect 413426 234498 413662 234734
rect 413106 234178 413342 234414
rect 413426 234178 413662 234414
rect 413106 198498 413342 198734
rect 413426 198498 413662 198734
rect 413106 198178 413342 198414
rect 413426 198178 413662 198414
rect 413106 162498 413342 162734
rect 413426 162498 413662 162734
rect 413106 162178 413342 162414
rect 413426 162178 413662 162414
rect 416826 709402 417062 709638
rect 417146 709402 417382 709638
rect 416826 709082 417062 709318
rect 417146 709082 417382 709318
rect 416826 670218 417062 670454
rect 417146 670218 417382 670454
rect 416826 669898 417062 670134
rect 417146 669898 417382 670134
rect 416826 634218 417062 634454
rect 417146 634218 417382 634454
rect 416826 633898 417062 634134
rect 417146 633898 417382 634134
rect 416826 598218 417062 598454
rect 417146 598218 417382 598454
rect 416826 597898 417062 598134
rect 417146 597898 417382 598134
rect 416826 562218 417062 562454
rect 417146 562218 417382 562454
rect 416826 561898 417062 562134
rect 417146 561898 417382 562134
rect 416826 526218 417062 526454
rect 417146 526218 417382 526454
rect 416826 525898 417062 526134
rect 417146 525898 417382 526134
rect 416826 490218 417062 490454
rect 417146 490218 417382 490454
rect 416826 489898 417062 490134
rect 417146 489898 417382 490134
rect 416826 454218 417062 454454
rect 417146 454218 417382 454454
rect 416826 453898 417062 454134
rect 417146 453898 417382 454134
rect 416826 418218 417062 418454
rect 417146 418218 417382 418454
rect 416826 417898 417062 418134
rect 417146 417898 417382 418134
rect 416826 382218 417062 382454
rect 417146 382218 417382 382454
rect 416826 381898 417062 382134
rect 417146 381898 417382 382134
rect 416826 346218 417062 346454
rect 417146 346218 417382 346454
rect 416826 345898 417062 346134
rect 417146 345898 417382 346134
rect 416826 310218 417062 310454
rect 417146 310218 417382 310454
rect 416826 309898 417062 310134
rect 417146 309898 417382 310134
rect 416826 274218 417062 274454
rect 417146 274218 417382 274454
rect 416826 273898 417062 274134
rect 417146 273898 417382 274134
rect 416826 238218 417062 238454
rect 417146 238218 417382 238454
rect 416826 237898 417062 238134
rect 417146 237898 417382 238134
rect 416826 202218 417062 202454
rect 417146 202218 417382 202454
rect 416826 201898 417062 202134
rect 417146 201898 417382 202134
rect 416826 166218 417062 166454
rect 417146 166218 417382 166454
rect 416826 165898 417062 166134
rect 417146 165898 417382 166134
rect 420546 710362 420782 710598
rect 420866 710362 421102 710598
rect 420546 710042 420782 710278
rect 420866 710042 421102 710278
rect 420546 673938 420782 674174
rect 420866 673938 421102 674174
rect 420546 673618 420782 673854
rect 420866 673618 421102 673854
rect 420546 637938 420782 638174
rect 420866 637938 421102 638174
rect 420546 637618 420782 637854
rect 420866 637618 421102 637854
rect 420546 601938 420782 602174
rect 420866 601938 421102 602174
rect 420546 601618 420782 601854
rect 420866 601618 421102 601854
rect 420546 565938 420782 566174
rect 420866 565938 421102 566174
rect 420546 565618 420782 565854
rect 420866 565618 421102 565854
rect 420546 529938 420782 530174
rect 420866 529938 421102 530174
rect 420546 529618 420782 529854
rect 420866 529618 421102 529854
rect 420546 493938 420782 494174
rect 420866 493938 421102 494174
rect 420546 493618 420782 493854
rect 420866 493618 421102 493854
rect 420546 457938 420782 458174
rect 420866 457938 421102 458174
rect 420546 457618 420782 457854
rect 420866 457618 421102 457854
rect 420546 421938 420782 422174
rect 420866 421938 421102 422174
rect 420546 421618 420782 421854
rect 420866 421618 421102 421854
rect 420546 385938 420782 386174
rect 420866 385938 421102 386174
rect 420546 385618 420782 385854
rect 420866 385618 421102 385854
rect 420546 349938 420782 350174
rect 420866 349938 421102 350174
rect 420546 349618 420782 349854
rect 420866 349618 421102 349854
rect 420546 313938 420782 314174
rect 420866 313938 421102 314174
rect 420546 313618 420782 313854
rect 420866 313618 421102 313854
rect 420546 277938 420782 278174
rect 420866 277938 421102 278174
rect 420546 277618 420782 277854
rect 420866 277618 421102 277854
rect 420546 241938 420782 242174
rect 420866 241938 421102 242174
rect 420546 241618 420782 241854
rect 420866 241618 421102 241854
rect 420546 205938 420782 206174
rect 420866 205938 421102 206174
rect 420546 205618 420782 205854
rect 420866 205618 421102 205854
rect 420546 169938 420782 170174
rect 420866 169938 421102 170174
rect 420546 169618 420782 169854
rect 420866 169618 421102 169854
rect 420546 133938 420782 134174
rect 420866 133938 421102 134174
rect 420546 133618 420782 133854
rect 420866 133618 421102 133854
rect 424266 711322 424502 711558
rect 424586 711322 424822 711558
rect 424266 711002 424502 711238
rect 424586 711002 424822 711238
rect 424266 677658 424502 677894
rect 424586 677658 424822 677894
rect 424266 677338 424502 677574
rect 424586 677338 424822 677574
rect 424266 641658 424502 641894
rect 424586 641658 424822 641894
rect 424266 641338 424502 641574
rect 424586 641338 424822 641574
rect 424266 605658 424502 605894
rect 424586 605658 424822 605894
rect 424266 605338 424502 605574
rect 424586 605338 424822 605574
rect 424266 569658 424502 569894
rect 424586 569658 424822 569894
rect 424266 569338 424502 569574
rect 424586 569338 424822 569574
rect 424266 533658 424502 533894
rect 424586 533658 424822 533894
rect 424266 533338 424502 533574
rect 424586 533338 424822 533574
rect 424266 497658 424502 497894
rect 424586 497658 424822 497894
rect 424266 497338 424502 497574
rect 424586 497338 424822 497574
rect 424266 461658 424502 461894
rect 424586 461658 424822 461894
rect 424266 461338 424502 461574
rect 424586 461338 424822 461574
rect 424266 425658 424502 425894
rect 424586 425658 424822 425894
rect 424266 425338 424502 425574
rect 424586 425338 424822 425574
rect 424266 389658 424502 389894
rect 424586 389658 424822 389894
rect 424266 389338 424502 389574
rect 424586 389338 424822 389574
rect 424266 353658 424502 353894
rect 424586 353658 424822 353894
rect 424266 353338 424502 353574
rect 424586 353338 424822 353574
rect 424266 317658 424502 317894
rect 424586 317658 424822 317894
rect 424266 317338 424502 317574
rect 424586 317338 424822 317574
rect 424266 281658 424502 281894
rect 424586 281658 424822 281894
rect 424266 281338 424502 281574
rect 424586 281338 424822 281574
rect 424266 245658 424502 245894
rect 424586 245658 424822 245894
rect 424266 245338 424502 245574
rect 424586 245338 424822 245574
rect 424266 209658 424502 209894
rect 424586 209658 424822 209894
rect 424266 209338 424502 209574
rect 424586 209338 424822 209574
rect 424266 173658 424502 173894
rect 424586 173658 424822 173894
rect 424266 173338 424502 173574
rect 424586 173338 424822 173574
rect 424266 137658 424502 137894
rect 424586 137658 424822 137894
rect 424266 137338 424502 137574
rect 424586 137338 424822 137574
rect 434226 704602 434462 704838
rect 434546 704602 434782 704838
rect 434226 704282 434462 704518
rect 434546 704282 434782 704518
rect 434226 687618 434462 687854
rect 434546 687618 434782 687854
rect 434226 687298 434462 687534
rect 434546 687298 434782 687534
rect 434226 651618 434462 651854
rect 434546 651618 434782 651854
rect 434226 651298 434462 651534
rect 434546 651298 434782 651534
rect 434226 615618 434462 615854
rect 434546 615618 434782 615854
rect 434226 615298 434462 615534
rect 434546 615298 434782 615534
rect 434226 579618 434462 579854
rect 434546 579618 434782 579854
rect 434226 579298 434462 579534
rect 434546 579298 434782 579534
rect 434226 543618 434462 543854
rect 434546 543618 434782 543854
rect 434226 543298 434462 543534
rect 434546 543298 434782 543534
rect 434226 507618 434462 507854
rect 434546 507618 434782 507854
rect 434226 507298 434462 507534
rect 434546 507298 434782 507534
rect 434226 471618 434462 471854
rect 434546 471618 434782 471854
rect 434226 471298 434462 471534
rect 434546 471298 434782 471534
rect 434226 435618 434462 435854
rect 434546 435618 434782 435854
rect 434226 435298 434462 435534
rect 434546 435298 434782 435534
rect 434226 399618 434462 399854
rect 434546 399618 434782 399854
rect 434226 399298 434462 399534
rect 434546 399298 434782 399534
rect 434226 363618 434462 363854
rect 434546 363618 434782 363854
rect 434226 363298 434462 363534
rect 434546 363298 434782 363534
rect 434226 327618 434462 327854
rect 434546 327618 434782 327854
rect 434226 327298 434462 327534
rect 434546 327298 434782 327534
rect 434226 291618 434462 291854
rect 434546 291618 434782 291854
rect 434226 291298 434462 291534
rect 434546 291298 434782 291534
rect 434226 255618 434462 255854
rect 434546 255618 434782 255854
rect 434226 255298 434462 255534
rect 434546 255298 434782 255534
rect 434226 219618 434462 219854
rect 434546 219618 434782 219854
rect 434226 219298 434462 219534
rect 434546 219298 434782 219534
rect 434226 183618 434462 183854
rect 434546 183618 434782 183854
rect 434226 183298 434462 183534
rect 434546 183298 434782 183534
rect 434226 147618 434462 147854
rect 434546 147618 434782 147854
rect 434226 147298 434462 147534
rect 434546 147298 434782 147534
rect 437946 705562 438182 705798
rect 438266 705562 438502 705798
rect 437946 705242 438182 705478
rect 438266 705242 438502 705478
rect 437946 691338 438182 691574
rect 438266 691338 438502 691574
rect 437946 691018 438182 691254
rect 438266 691018 438502 691254
rect 437946 655338 438182 655574
rect 438266 655338 438502 655574
rect 437946 655018 438182 655254
rect 438266 655018 438502 655254
rect 437946 619338 438182 619574
rect 438266 619338 438502 619574
rect 437946 619018 438182 619254
rect 438266 619018 438502 619254
rect 437946 583338 438182 583574
rect 438266 583338 438502 583574
rect 437946 583018 438182 583254
rect 438266 583018 438502 583254
rect 437946 547338 438182 547574
rect 438266 547338 438502 547574
rect 437946 547018 438182 547254
rect 438266 547018 438502 547254
rect 437946 511338 438182 511574
rect 438266 511338 438502 511574
rect 437946 511018 438182 511254
rect 438266 511018 438502 511254
rect 437946 475338 438182 475574
rect 438266 475338 438502 475574
rect 437946 475018 438182 475254
rect 438266 475018 438502 475254
rect 437946 439338 438182 439574
rect 438266 439338 438502 439574
rect 437946 439018 438182 439254
rect 438266 439018 438502 439254
rect 437946 403338 438182 403574
rect 438266 403338 438502 403574
rect 437946 403018 438182 403254
rect 438266 403018 438502 403254
rect 437946 367338 438182 367574
rect 438266 367338 438502 367574
rect 437946 367018 438182 367254
rect 438266 367018 438502 367254
rect 437946 331338 438182 331574
rect 438266 331338 438502 331574
rect 437946 331018 438182 331254
rect 438266 331018 438502 331254
rect 437946 295338 438182 295574
rect 438266 295338 438502 295574
rect 437946 295018 438182 295254
rect 438266 295018 438502 295254
rect 437946 259338 438182 259574
rect 438266 259338 438502 259574
rect 437946 259018 438182 259254
rect 438266 259018 438502 259254
rect 437946 223338 438182 223574
rect 438266 223338 438502 223574
rect 437946 223018 438182 223254
rect 438266 223018 438502 223254
rect 437946 187338 438182 187574
rect 438266 187338 438502 187574
rect 437946 187018 438182 187254
rect 438266 187018 438502 187254
rect 437946 151338 438182 151574
rect 438266 151338 438502 151574
rect 437946 151018 438182 151254
rect 438266 151018 438502 151254
rect 441666 706522 441902 706758
rect 441986 706522 442222 706758
rect 441666 706202 441902 706438
rect 441986 706202 442222 706438
rect 441666 695058 441902 695294
rect 441986 695058 442222 695294
rect 441666 694738 441902 694974
rect 441986 694738 442222 694974
rect 441666 659058 441902 659294
rect 441986 659058 442222 659294
rect 441666 658738 441902 658974
rect 441986 658738 442222 658974
rect 441666 623058 441902 623294
rect 441986 623058 442222 623294
rect 441666 622738 441902 622974
rect 441986 622738 442222 622974
rect 441666 587058 441902 587294
rect 441986 587058 442222 587294
rect 441666 586738 441902 586974
rect 441986 586738 442222 586974
rect 441666 551058 441902 551294
rect 441986 551058 442222 551294
rect 441666 550738 441902 550974
rect 441986 550738 442222 550974
rect 441666 515058 441902 515294
rect 441986 515058 442222 515294
rect 441666 514738 441902 514974
rect 441986 514738 442222 514974
rect 441666 479058 441902 479294
rect 441986 479058 442222 479294
rect 441666 478738 441902 478974
rect 441986 478738 442222 478974
rect 441666 443058 441902 443294
rect 441986 443058 442222 443294
rect 441666 442738 441902 442974
rect 441986 442738 442222 442974
rect 441666 407058 441902 407294
rect 441986 407058 442222 407294
rect 441666 406738 441902 406974
rect 441986 406738 442222 406974
rect 441666 371058 441902 371294
rect 441986 371058 442222 371294
rect 441666 370738 441902 370974
rect 441986 370738 442222 370974
rect 441666 335058 441902 335294
rect 441986 335058 442222 335294
rect 441666 334738 441902 334974
rect 441986 334738 442222 334974
rect 441666 299058 441902 299294
rect 441986 299058 442222 299294
rect 441666 298738 441902 298974
rect 441986 298738 442222 298974
rect 441666 263058 441902 263294
rect 441986 263058 442222 263294
rect 441666 262738 441902 262974
rect 441986 262738 442222 262974
rect 441666 227058 441902 227294
rect 441986 227058 442222 227294
rect 441666 226738 441902 226974
rect 441986 226738 442222 226974
rect 441666 191058 441902 191294
rect 441986 191058 442222 191294
rect 441666 190738 441902 190974
rect 441986 190738 442222 190974
rect 441666 155058 441902 155294
rect 441986 155058 442222 155294
rect 441666 154738 441902 154974
rect 441986 154738 442222 154974
rect 445386 707482 445622 707718
rect 445706 707482 445942 707718
rect 445386 707162 445622 707398
rect 445706 707162 445942 707398
rect 445386 698778 445622 699014
rect 445706 698778 445942 699014
rect 445386 698458 445622 698694
rect 445706 698458 445942 698694
rect 445386 662778 445622 663014
rect 445706 662778 445942 663014
rect 445386 662458 445622 662694
rect 445706 662458 445942 662694
rect 445386 626778 445622 627014
rect 445706 626778 445942 627014
rect 445386 626458 445622 626694
rect 445706 626458 445942 626694
rect 445386 590778 445622 591014
rect 445706 590778 445942 591014
rect 445386 590458 445622 590694
rect 445706 590458 445942 590694
rect 445386 554778 445622 555014
rect 445706 554778 445942 555014
rect 445386 554458 445622 554694
rect 445706 554458 445942 554694
rect 445386 518778 445622 519014
rect 445706 518778 445942 519014
rect 445386 518458 445622 518694
rect 445706 518458 445942 518694
rect 445386 482778 445622 483014
rect 445706 482778 445942 483014
rect 445386 482458 445622 482694
rect 445706 482458 445942 482694
rect 445386 446778 445622 447014
rect 445706 446778 445942 447014
rect 445386 446458 445622 446694
rect 445706 446458 445942 446694
rect 445386 410778 445622 411014
rect 445706 410778 445942 411014
rect 445386 410458 445622 410694
rect 445706 410458 445942 410694
rect 445386 374778 445622 375014
rect 445706 374778 445942 375014
rect 445386 374458 445622 374694
rect 445706 374458 445942 374694
rect 445386 338778 445622 339014
rect 445706 338778 445942 339014
rect 445386 338458 445622 338694
rect 445706 338458 445942 338694
rect 445386 302778 445622 303014
rect 445706 302778 445942 303014
rect 445386 302458 445622 302694
rect 445706 302458 445942 302694
rect 445386 266778 445622 267014
rect 445706 266778 445942 267014
rect 445386 266458 445622 266694
rect 445706 266458 445942 266694
rect 445386 230778 445622 231014
rect 445706 230778 445942 231014
rect 445386 230458 445622 230694
rect 445706 230458 445942 230694
rect 445386 194778 445622 195014
rect 445706 194778 445942 195014
rect 445386 194458 445622 194694
rect 445706 194458 445942 194694
rect 445386 158778 445622 159014
rect 445706 158778 445942 159014
rect 445386 158458 445622 158694
rect 445706 158458 445942 158694
rect 449106 708442 449342 708678
rect 449426 708442 449662 708678
rect 449106 708122 449342 708358
rect 449426 708122 449662 708358
rect 449106 666498 449342 666734
rect 449426 666498 449662 666734
rect 449106 666178 449342 666414
rect 449426 666178 449662 666414
rect 449106 630498 449342 630734
rect 449426 630498 449662 630734
rect 449106 630178 449342 630414
rect 449426 630178 449662 630414
rect 449106 594498 449342 594734
rect 449426 594498 449662 594734
rect 449106 594178 449342 594414
rect 449426 594178 449662 594414
rect 449106 558498 449342 558734
rect 449426 558498 449662 558734
rect 449106 558178 449342 558414
rect 449426 558178 449662 558414
rect 449106 522498 449342 522734
rect 449426 522498 449662 522734
rect 449106 522178 449342 522414
rect 449426 522178 449662 522414
rect 449106 486498 449342 486734
rect 449426 486498 449662 486734
rect 449106 486178 449342 486414
rect 449426 486178 449662 486414
rect 449106 450498 449342 450734
rect 449426 450498 449662 450734
rect 449106 450178 449342 450414
rect 449426 450178 449662 450414
rect 449106 414498 449342 414734
rect 449426 414498 449662 414734
rect 449106 414178 449342 414414
rect 449426 414178 449662 414414
rect 449106 378498 449342 378734
rect 449426 378498 449662 378734
rect 449106 378178 449342 378414
rect 449426 378178 449662 378414
rect 449106 342498 449342 342734
rect 449426 342498 449662 342734
rect 449106 342178 449342 342414
rect 449426 342178 449662 342414
rect 449106 306498 449342 306734
rect 449426 306498 449662 306734
rect 449106 306178 449342 306414
rect 449426 306178 449662 306414
rect 449106 270498 449342 270734
rect 449426 270498 449662 270734
rect 449106 270178 449342 270414
rect 449426 270178 449662 270414
rect 449106 234498 449342 234734
rect 449426 234498 449662 234734
rect 449106 234178 449342 234414
rect 449426 234178 449662 234414
rect 449106 198498 449342 198734
rect 449426 198498 449662 198734
rect 449106 198178 449342 198414
rect 449426 198178 449662 198414
rect 449106 162498 449342 162734
rect 449426 162498 449662 162734
rect 449106 162178 449342 162414
rect 449426 162178 449662 162414
rect 452826 709402 453062 709638
rect 453146 709402 453382 709638
rect 452826 709082 453062 709318
rect 453146 709082 453382 709318
rect 452826 670218 453062 670454
rect 453146 670218 453382 670454
rect 452826 669898 453062 670134
rect 453146 669898 453382 670134
rect 452826 634218 453062 634454
rect 453146 634218 453382 634454
rect 452826 633898 453062 634134
rect 453146 633898 453382 634134
rect 452826 598218 453062 598454
rect 453146 598218 453382 598454
rect 452826 597898 453062 598134
rect 453146 597898 453382 598134
rect 452826 562218 453062 562454
rect 453146 562218 453382 562454
rect 452826 561898 453062 562134
rect 453146 561898 453382 562134
rect 452826 526218 453062 526454
rect 453146 526218 453382 526454
rect 452826 525898 453062 526134
rect 453146 525898 453382 526134
rect 452826 490218 453062 490454
rect 453146 490218 453382 490454
rect 452826 489898 453062 490134
rect 453146 489898 453382 490134
rect 452826 454218 453062 454454
rect 453146 454218 453382 454454
rect 452826 453898 453062 454134
rect 453146 453898 453382 454134
rect 452826 418218 453062 418454
rect 453146 418218 453382 418454
rect 452826 417898 453062 418134
rect 453146 417898 453382 418134
rect 452826 382218 453062 382454
rect 453146 382218 453382 382454
rect 452826 381898 453062 382134
rect 453146 381898 453382 382134
rect 452826 346218 453062 346454
rect 453146 346218 453382 346454
rect 452826 345898 453062 346134
rect 453146 345898 453382 346134
rect 452826 310218 453062 310454
rect 453146 310218 453382 310454
rect 452826 309898 453062 310134
rect 453146 309898 453382 310134
rect 452826 274218 453062 274454
rect 453146 274218 453382 274454
rect 452826 273898 453062 274134
rect 453146 273898 453382 274134
rect 452826 238218 453062 238454
rect 453146 238218 453382 238454
rect 452826 237898 453062 238134
rect 453146 237898 453382 238134
rect 452826 202218 453062 202454
rect 453146 202218 453382 202454
rect 452826 201898 453062 202134
rect 453146 201898 453382 202134
rect 452826 166218 453062 166454
rect 453146 166218 453382 166454
rect 452826 165898 453062 166134
rect 453146 165898 453382 166134
rect 409386 122778 409622 123014
rect 409706 122778 409942 123014
rect 409386 122458 409622 122694
rect 409706 122458 409942 122694
rect 452826 130218 453062 130454
rect 453146 130218 453382 130454
rect 452826 129898 453062 130134
rect 453146 129898 453382 130134
rect 419610 115338 419846 115574
rect 419610 115018 419846 115254
rect 450330 115338 450566 115574
rect 450330 115018 450566 115254
rect 434970 111618 435206 111854
rect 434970 111298 435206 111534
rect 409386 86778 409622 87014
rect 409706 86778 409942 87014
rect 409386 86458 409622 86694
rect 409706 86458 409942 86694
rect 405666 47058 405902 47294
rect 405986 47058 406222 47294
rect 405666 46738 405902 46974
rect 405986 46738 406222 46974
rect 405666 11058 405902 11294
rect 405986 11058 406222 11294
rect 405666 10738 405902 10974
rect 405986 10738 406222 10974
rect 452826 94218 453062 94454
rect 453146 94218 453382 94454
rect 452826 93898 453062 94134
rect 453146 93898 453382 94134
rect 409386 50778 409622 51014
rect 409706 50778 409942 51014
rect 409386 50458 409622 50694
rect 409706 50458 409942 50694
rect 409386 14778 409622 15014
rect 409706 14778 409942 15014
rect 409386 14458 409622 14694
rect 409706 14458 409942 14694
rect 405666 -2502 405902 -2266
rect 405986 -2502 406222 -2266
rect 405666 -2822 405902 -2586
rect 405986 -2822 406222 -2586
rect 413106 54498 413342 54734
rect 413426 54498 413662 54734
rect 413106 54178 413342 54414
rect 413426 54178 413662 54414
rect 413106 18498 413342 18734
rect 413426 18498 413662 18734
rect 413106 18178 413342 18414
rect 413426 18178 413662 18414
rect 409386 -3462 409622 -3226
rect 409706 -3462 409942 -3226
rect 409386 -3782 409622 -3546
rect 409706 -3782 409942 -3546
rect 413106 -4422 413342 -4186
rect 413426 -4422 413662 -4186
rect 413106 -4742 413342 -4506
rect 413426 -4742 413662 -4506
rect 416826 58218 417062 58454
rect 417146 58218 417382 58454
rect 416826 57898 417062 58134
rect 417146 57898 417382 58134
rect 416826 22218 417062 22454
rect 417146 22218 417382 22454
rect 416826 21898 417062 22134
rect 417146 21898 417382 22134
rect 416826 -5382 417062 -5146
rect 417146 -5382 417382 -5146
rect 416826 -5702 417062 -5466
rect 417146 -5702 417382 -5466
rect 420546 61938 420782 62174
rect 420866 61938 421102 62174
rect 420546 61618 420782 61854
rect 420866 61618 421102 61854
rect 420546 25938 420782 26174
rect 420866 25938 421102 26174
rect 420546 25618 420782 25854
rect 420866 25618 421102 25854
rect 420546 -6342 420782 -6106
rect 420866 -6342 421102 -6106
rect 420546 -6662 420782 -6426
rect 420866 -6662 421102 -6426
rect 424266 65658 424502 65894
rect 424586 65658 424822 65894
rect 424266 65338 424502 65574
rect 424586 65338 424822 65574
rect 424266 29658 424502 29894
rect 424586 29658 424822 29894
rect 424266 29338 424502 29574
rect 424586 29338 424822 29574
rect 434226 75618 434462 75854
rect 434546 75618 434782 75854
rect 434226 75298 434462 75534
rect 434546 75298 434782 75534
rect 434226 39618 434462 39854
rect 434546 39618 434782 39854
rect 434226 39298 434462 39534
rect 434546 39298 434782 39534
rect 431638 9062 431874 9298
rect 424266 -7302 424502 -7066
rect 424586 -7302 424822 -7066
rect 424266 -7622 424502 -7386
rect 424586 -7622 424822 -7386
rect 434226 3618 434462 3854
rect 434546 3618 434782 3854
rect 434226 3298 434462 3534
rect 434546 3298 434782 3534
rect 434226 -582 434462 -346
rect 434546 -582 434782 -346
rect 434226 -902 434462 -666
rect 434546 -902 434782 -666
rect 437946 79338 438182 79574
rect 438266 79338 438502 79574
rect 437946 79018 438182 79254
rect 438266 79018 438502 79254
rect 437946 43338 438182 43574
rect 438266 43338 438502 43574
rect 437946 43018 438182 43254
rect 438266 43018 438502 43254
rect 437946 7338 438182 7574
rect 438266 7338 438502 7574
rect 437946 7018 438182 7254
rect 438266 7018 438502 7254
rect 437946 -1542 438182 -1306
rect 438266 -1542 438502 -1306
rect 437946 -1862 438182 -1626
rect 438266 -1862 438502 -1626
rect 441666 47058 441902 47294
rect 441986 47058 442222 47294
rect 441666 46738 441902 46974
rect 441986 46738 442222 46974
rect 441666 11058 441902 11294
rect 441986 11058 442222 11294
rect 441666 10738 441902 10974
rect 441986 10738 442222 10974
rect 441666 -2502 441902 -2266
rect 441986 -2502 442222 -2266
rect 441666 -2822 441902 -2586
rect 441986 -2822 442222 -2586
rect 445386 50778 445622 51014
rect 445706 50778 445942 51014
rect 445386 50458 445622 50694
rect 445706 50458 445942 50694
rect 445386 14778 445622 15014
rect 445706 14778 445942 15014
rect 445386 14458 445622 14694
rect 445706 14458 445942 14694
rect 445386 -3462 445622 -3226
rect 445706 -3462 445942 -3226
rect 445386 -3782 445622 -3546
rect 445706 -3782 445942 -3546
rect 449106 54498 449342 54734
rect 449426 54498 449662 54734
rect 449106 54178 449342 54414
rect 449426 54178 449662 54414
rect 449106 18498 449342 18734
rect 449426 18498 449662 18734
rect 449106 18178 449342 18414
rect 449426 18178 449662 18414
rect 449106 -4422 449342 -4186
rect 449426 -4422 449662 -4186
rect 449106 -4742 449342 -4506
rect 449426 -4742 449662 -4506
rect 452826 58218 453062 58454
rect 453146 58218 453382 58454
rect 452826 57898 453062 58134
rect 453146 57898 453382 58134
rect 452826 22218 453062 22454
rect 453146 22218 453382 22454
rect 452826 21898 453062 22134
rect 453146 21898 453382 22134
rect 452826 -5382 453062 -5146
rect 453146 -5382 453382 -5146
rect 452826 -5702 453062 -5466
rect 453146 -5702 453382 -5466
rect 456546 710362 456782 710598
rect 456866 710362 457102 710598
rect 456546 710042 456782 710278
rect 456866 710042 457102 710278
rect 456546 673938 456782 674174
rect 456866 673938 457102 674174
rect 456546 673618 456782 673854
rect 456866 673618 457102 673854
rect 456546 637938 456782 638174
rect 456866 637938 457102 638174
rect 456546 637618 456782 637854
rect 456866 637618 457102 637854
rect 456546 601938 456782 602174
rect 456866 601938 457102 602174
rect 456546 601618 456782 601854
rect 456866 601618 457102 601854
rect 456546 565938 456782 566174
rect 456866 565938 457102 566174
rect 456546 565618 456782 565854
rect 456866 565618 457102 565854
rect 456546 529938 456782 530174
rect 456866 529938 457102 530174
rect 456546 529618 456782 529854
rect 456866 529618 457102 529854
rect 456546 493938 456782 494174
rect 456866 493938 457102 494174
rect 456546 493618 456782 493854
rect 456866 493618 457102 493854
rect 456546 457938 456782 458174
rect 456866 457938 457102 458174
rect 456546 457618 456782 457854
rect 456866 457618 457102 457854
rect 456546 421938 456782 422174
rect 456866 421938 457102 422174
rect 456546 421618 456782 421854
rect 456866 421618 457102 421854
rect 456546 385938 456782 386174
rect 456866 385938 457102 386174
rect 456546 385618 456782 385854
rect 456866 385618 457102 385854
rect 456546 349938 456782 350174
rect 456866 349938 457102 350174
rect 456546 349618 456782 349854
rect 456866 349618 457102 349854
rect 456546 313938 456782 314174
rect 456866 313938 457102 314174
rect 456546 313618 456782 313854
rect 456866 313618 457102 313854
rect 456546 277938 456782 278174
rect 456866 277938 457102 278174
rect 456546 277618 456782 277854
rect 456866 277618 457102 277854
rect 456546 241938 456782 242174
rect 456866 241938 457102 242174
rect 456546 241618 456782 241854
rect 456866 241618 457102 241854
rect 456546 205938 456782 206174
rect 456866 205938 457102 206174
rect 456546 205618 456782 205854
rect 456866 205618 457102 205854
rect 456546 169938 456782 170174
rect 456866 169938 457102 170174
rect 456546 169618 456782 169854
rect 456866 169618 457102 169854
rect 456546 133938 456782 134174
rect 456866 133938 457102 134174
rect 456546 133618 456782 133854
rect 456866 133618 457102 133854
rect 456546 97938 456782 98174
rect 456866 97938 457102 98174
rect 456546 97618 456782 97854
rect 456866 97618 457102 97854
rect 456546 61938 456782 62174
rect 456866 61938 457102 62174
rect 456546 61618 456782 61854
rect 456866 61618 457102 61854
rect 456546 25938 456782 26174
rect 456866 25938 457102 26174
rect 456546 25618 456782 25854
rect 456866 25618 457102 25854
rect 456546 -6342 456782 -6106
rect 456866 -6342 457102 -6106
rect 456546 -6662 456782 -6426
rect 456866 -6662 457102 -6426
rect 460266 711322 460502 711558
rect 460586 711322 460822 711558
rect 460266 711002 460502 711238
rect 460586 711002 460822 711238
rect 460266 677658 460502 677894
rect 460586 677658 460822 677894
rect 460266 677338 460502 677574
rect 460586 677338 460822 677574
rect 460266 641658 460502 641894
rect 460586 641658 460822 641894
rect 460266 641338 460502 641574
rect 460586 641338 460822 641574
rect 460266 605658 460502 605894
rect 460586 605658 460822 605894
rect 460266 605338 460502 605574
rect 460586 605338 460822 605574
rect 460266 569658 460502 569894
rect 460586 569658 460822 569894
rect 460266 569338 460502 569574
rect 460586 569338 460822 569574
rect 460266 533658 460502 533894
rect 460586 533658 460822 533894
rect 460266 533338 460502 533574
rect 460586 533338 460822 533574
rect 460266 497658 460502 497894
rect 460586 497658 460822 497894
rect 460266 497338 460502 497574
rect 460586 497338 460822 497574
rect 460266 461658 460502 461894
rect 460586 461658 460822 461894
rect 460266 461338 460502 461574
rect 460586 461338 460822 461574
rect 460266 425658 460502 425894
rect 460586 425658 460822 425894
rect 460266 425338 460502 425574
rect 460586 425338 460822 425574
rect 460266 389658 460502 389894
rect 460586 389658 460822 389894
rect 460266 389338 460502 389574
rect 460586 389338 460822 389574
rect 460266 353658 460502 353894
rect 460586 353658 460822 353894
rect 460266 353338 460502 353574
rect 460586 353338 460822 353574
rect 460266 317658 460502 317894
rect 460586 317658 460822 317894
rect 460266 317338 460502 317574
rect 460586 317338 460822 317574
rect 460266 281658 460502 281894
rect 460586 281658 460822 281894
rect 460266 281338 460502 281574
rect 460586 281338 460822 281574
rect 460266 245658 460502 245894
rect 460586 245658 460822 245894
rect 460266 245338 460502 245574
rect 460586 245338 460822 245574
rect 460266 209658 460502 209894
rect 460586 209658 460822 209894
rect 460266 209338 460502 209574
rect 460586 209338 460822 209574
rect 460266 173658 460502 173894
rect 460586 173658 460822 173894
rect 460266 173338 460502 173574
rect 460586 173338 460822 173574
rect 460266 137658 460502 137894
rect 460586 137658 460822 137894
rect 460266 137338 460502 137574
rect 460586 137338 460822 137574
rect 460266 101658 460502 101894
rect 460586 101658 460822 101894
rect 460266 101338 460502 101574
rect 460586 101338 460822 101574
rect 460266 65658 460502 65894
rect 460586 65658 460822 65894
rect 460266 65338 460502 65574
rect 460586 65338 460822 65574
rect 460266 29658 460502 29894
rect 460586 29658 460822 29894
rect 460266 29338 460502 29574
rect 460586 29338 460822 29574
rect 460266 -7302 460502 -7066
rect 460586 -7302 460822 -7066
rect 460266 -7622 460502 -7386
rect 460586 -7622 460822 -7386
rect 470226 704602 470462 704838
rect 470546 704602 470782 704838
rect 470226 704282 470462 704518
rect 470546 704282 470782 704518
rect 470226 687618 470462 687854
rect 470546 687618 470782 687854
rect 470226 687298 470462 687534
rect 470546 687298 470782 687534
rect 470226 651618 470462 651854
rect 470546 651618 470782 651854
rect 470226 651298 470462 651534
rect 470546 651298 470782 651534
rect 470226 615618 470462 615854
rect 470546 615618 470782 615854
rect 470226 615298 470462 615534
rect 470546 615298 470782 615534
rect 470226 579618 470462 579854
rect 470546 579618 470782 579854
rect 470226 579298 470462 579534
rect 470546 579298 470782 579534
rect 470226 543618 470462 543854
rect 470546 543618 470782 543854
rect 470226 543298 470462 543534
rect 470546 543298 470782 543534
rect 470226 507618 470462 507854
rect 470546 507618 470782 507854
rect 470226 507298 470462 507534
rect 470546 507298 470782 507534
rect 470226 471618 470462 471854
rect 470546 471618 470782 471854
rect 470226 471298 470462 471534
rect 470546 471298 470782 471534
rect 470226 435618 470462 435854
rect 470546 435618 470782 435854
rect 470226 435298 470462 435534
rect 470546 435298 470782 435534
rect 470226 399618 470462 399854
rect 470546 399618 470782 399854
rect 470226 399298 470462 399534
rect 470546 399298 470782 399534
rect 470226 363618 470462 363854
rect 470546 363618 470782 363854
rect 470226 363298 470462 363534
rect 470546 363298 470782 363534
rect 470226 327618 470462 327854
rect 470546 327618 470782 327854
rect 470226 327298 470462 327534
rect 470546 327298 470782 327534
rect 470226 291618 470462 291854
rect 470546 291618 470782 291854
rect 470226 291298 470462 291534
rect 470546 291298 470782 291534
rect 470226 255618 470462 255854
rect 470546 255618 470782 255854
rect 470226 255298 470462 255534
rect 470546 255298 470782 255534
rect 470226 219618 470462 219854
rect 470546 219618 470782 219854
rect 470226 219298 470462 219534
rect 470546 219298 470782 219534
rect 470226 183618 470462 183854
rect 470546 183618 470782 183854
rect 470226 183298 470462 183534
rect 470546 183298 470782 183534
rect 470226 147618 470462 147854
rect 470546 147618 470782 147854
rect 470226 147298 470462 147534
rect 470546 147298 470782 147534
rect 470226 111618 470462 111854
rect 470546 111618 470782 111854
rect 470226 111298 470462 111534
rect 470546 111298 470782 111534
rect 470226 75618 470462 75854
rect 470546 75618 470782 75854
rect 470226 75298 470462 75534
rect 470546 75298 470782 75534
rect 470226 39618 470462 39854
rect 470546 39618 470782 39854
rect 470226 39298 470462 39534
rect 470546 39298 470782 39534
rect 470226 3618 470462 3854
rect 470546 3618 470782 3854
rect 470226 3298 470462 3534
rect 470546 3298 470782 3534
rect 470226 -582 470462 -346
rect 470546 -582 470782 -346
rect 470226 -902 470462 -666
rect 470546 -902 470782 -666
rect 473946 705562 474182 705798
rect 474266 705562 474502 705798
rect 473946 705242 474182 705478
rect 474266 705242 474502 705478
rect 473946 691338 474182 691574
rect 474266 691338 474502 691574
rect 473946 691018 474182 691254
rect 474266 691018 474502 691254
rect 473946 655338 474182 655574
rect 474266 655338 474502 655574
rect 473946 655018 474182 655254
rect 474266 655018 474502 655254
rect 473946 619338 474182 619574
rect 474266 619338 474502 619574
rect 473946 619018 474182 619254
rect 474266 619018 474502 619254
rect 473946 583338 474182 583574
rect 474266 583338 474502 583574
rect 473946 583018 474182 583254
rect 474266 583018 474502 583254
rect 473946 547338 474182 547574
rect 474266 547338 474502 547574
rect 473946 547018 474182 547254
rect 474266 547018 474502 547254
rect 473946 511338 474182 511574
rect 474266 511338 474502 511574
rect 473946 511018 474182 511254
rect 474266 511018 474502 511254
rect 473946 475338 474182 475574
rect 474266 475338 474502 475574
rect 473946 475018 474182 475254
rect 474266 475018 474502 475254
rect 473946 439338 474182 439574
rect 474266 439338 474502 439574
rect 473946 439018 474182 439254
rect 474266 439018 474502 439254
rect 473946 403338 474182 403574
rect 474266 403338 474502 403574
rect 473946 403018 474182 403254
rect 474266 403018 474502 403254
rect 473946 367338 474182 367574
rect 474266 367338 474502 367574
rect 473946 367018 474182 367254
rect 474266 367018 474502 367254
rect 473946 331338 474182 331574
rect 474266 331338 474502 331574
rect 473946 331018 474182 331254
rect 474266 331018 474502 331254
rect 473946 295338 474182 295574
rect 474266 295338 474502 295574
rect 473946 295018 474182 295254
rect 474266 295018 474502 295254
rect 473946 259338 474182 259574
rect 474266 259338 474502 259574
rect 473946 259018 474182 259254
rect 474266 259018 474502 259254
rect 473946 223338 474182 223574
rect 474266 223338 474502 223574
rect 473946 223018 474182 223254
rect 474266 223018 474502 223254
rect 473946 187338 474182 187574
rect 474266 187338 474502 187574
rect 473946 187018 474182 187254
rect 474266 187018 474502 187254
rect 473946 151338 474182 151574
rect 474266 151338 474502 151574
rect 473946 151018 474182 151254
rect 474266 151018 474502 151254
rect 473946 115338 474182 115574
rect 474266 115338 474502 115574
rect 473946 115018 474182 115254
rect 474266 115018 474502 115254
rect 473946 79338 474182 79574
rect 474266 79338 474502 79574
rect 473946 79018 474182 79254
rect 474266 79018 474502 79254
rect 473946 43338 474182 43574
rect 474266 43338 474502 43574
rect 473946 43018 474182 43254
rect 474266 43018 474502 43254
rect 473946 7338 474182 7574
rect 474266 7338 474502 7574
rect 473946 7018 474182 7254
rect 474266 7018 474502 7254
rect 473946 -1542 474182 -1306
rect 474266 -1542 474502 -1306
rect 473946 -1862 474182 -1626
rect 474266 -1862 474502 -1626
rect 477666 706522 477902 706758
rect 477986 706522 478222 706758
rect 477666 706202 477902 706438
rect 477986 706202 478222 706438
rect 477666 695058 477902 695294
rect 477986 695058 478222 695294
rect 477666 694738 477902 694974
rect 477986 694738 478222 694974
rect 477666 659058 477902 659294
rect 477986 659058 478222 659294
rect 477666 658738 477902 658974
rect 477986 658738 478222 658974
rect 477666 623058 477902 623294
rect 477986 623058 478222 623294
rect 477666 622738 477902 622974
rect 477986 622738 478222 622974
rect 477666 587058 477902 587294
rect 477986 587058 478222 587294
rect 477666 586738 477902 586974
rect 477986 586738 478222 586974
rect 477666 551058 477902 551294
rect 477986 551058 478222 551294
rect 477666 550738 477902 550974
rect 477986 550738 478222 550974
rect 477666 515058 477902 515294
rect 477986 515058 478222 515294
rect 477666 514738 477902 514974
rect 477986 514738 478222 514974
rect 477666 479058 477902 479294
rect 477986 479058 478222 479294
rect 477666 478738 477902 478974
rect 477986 478738 478222 478974
rect 477666 443058 477902 443294
rect 477986 443058 478222 443294
rect 477666 442738 477902 442974
rect 477986 442738 478222 442974
rect 477666 407058 477902 407294
rect 477986 407058 478222 407294
rect 477666 406738 477902 406974
rect 477986 406738 478222 406974
rect 477666 371058 477902 371294
rect 477986 371058 478222 371294
rect 477666 370738 477902 370974
rect 477986 370738 478222 370974
rect 477666 335058 477902 335294
rect 477986 335058 478222 335294
rect 477666 334738 477902 334974
rect 477986 334738 478222 334974
rect 477666 299058 477902 299294
rect 477986 299058 478222 299294
rect 477666 298738 477902 298974
rect 477986 298738 478222 298974
rect 477666 263058 477902 263294
rect 477986 263058 478222 263294
rect 477666 262738 477902 262974
rect 477986 262738 478222 262974
rect 477666 227058 477902 227294
rect 477986 227058 478222 227294
rect 477666 226738 477902 226974
rect 477986 226738 478222 226974
rect 477666 191058 477902 191294
rect 477986 191058 478222 191294
rect 477666 190738 477902 190974
rect 477986 190738 478222 190974
rect 477666 155058 477902 155294
rect 477986 155058 478222 155294
rect 477666 154738 477902 154974
rect 477986 154738 478222 154974
rect 477666 119058 477902 119294
rect 477986 119058 478222 119294
rect 477666 118738 477902 118974
rect 477986 118738 478222 118974
rect 477666 83058 477902 83294
rect 477986 83058 478222 83294
rect 477666 82738 477902 82974
rect 477986 82738 478222 82974
rect 477666 47058 477902 47294
rect 477986 47058 478222 47294
rect 477666 46738 477902 46974
rect 477986 46738 478222 46974
rect 477666 11058 477902 11294
rect 477986 11058 478222 11294
rect 477666 10738 477902 10974
rect 477986 10738 478222 10974
rect 477666 -2502 477902 -2266
rect 477986 -2502 478222 -2266
rect 477666 -2822 477902 -2586
rect 477986 -2822 478222 -2586
rect 481386 707482 481622 707718
rect 481706 707482 481942 707718
rect 481386 707162 481622 707398
rect 481706 707162 481942 707398
rect 481386 698778 481622 699014
rect 481706 698778 481942 699014
rect 481386 698458 481622 698694
rect 481706 698458 481942 698694
rect 481386 662778 481622 663014
rect 481706 662778 481942 663014
rect 481386 662458 481622 662694
rect 481706 662458 481942 662694
rect 481386 626778 481622 627014
rect 481706 626778 481942 627014
rect 481386 626458 481622 626694
rect 481706 626458 481942 626694
rect 481386 590778 481622 591014
rect 481706 590778 481942 591014
rect 481386 590458 481622 590694
rect 481706 590458 481942 590694
rect 481386 554778 481622 555014
rect 481706 554778 481942 555014
rect 481386 554458 481622 554694
rect 481706 554458 481942 554694
rect 481386 518778 481622 519014
rect 481706 518778 481942 519014
rect 481386 518458 481622 518694
rect 481706 518458 481942 518694
rect 481386 482778 481622 483014
rect 481706 482778 481942 483014
rect 481386 482458 481622 482694
rect 481706 482458 481942 482694
rect 481386 446778 481622 447014
rect 481706 446778 481942 447014
rect 481386 446458 481622 446694
rect 481706 446458 481942 446694
rect 481386 410778 481622 411014
rect 481706 410778 481942 411014
rect 481386 410458 481622 410694
rect 481706 410458 481942 410694
rect 481386 374778 481622 375014
rect 481706 374778 481942 375014
rect 481386 374458 481622 374694
rect 481706 374458 481942 374694
rect 481386 338778 481622 339014
rect 481706 338778 481942 339014
rect 481386 338458 481622 338694
rect 481706 338458 481942 338694
rect 481386 302778 481622 303014
rect 481706 302778 481942 303014
rect 481386 302458 481622 302694
rect 481706 302458 481942 302694
rect 481386 266778 481622 267014
rect 481706 266778 481942 267014
rect 481386 266458 481622 266694
rect 481706 266458 481942 266694
rect 481386 230778 481622 231014
rect 481706 230778 481942 231014
rect 481386 230458 481622 230694
rect 481706 230458 481942 230694
rect 481386 194778 481622 195014
rect 481706 194778 481942 195014
rect 481386 194458 481622 194694
rect 481706 194458 481942 194694
rect 481386 158778 481622 159014
rect 481706 158778 481942 159014
rect 481386 158458 481622 158694
rect 481706 158458 481942 158694
rect 481386 122778 481622 123014
rect 481706 122778 481942 123014
rect 481386 122458 481622 122694
rect 481706 122458 481942 122694
rect 481386 86778 481622 87014
rect 481706 86778 481942 87014
rect 481386 86458 481622 86694
rect 481706 86458 481942 86694
rect 481386 50778 481622 51014
rect 481706 50778 481942 51014
rect 481386 50458 481622 50694
rect 481706 50458 481942 50694
rect 481386 14778 481622 15014
rect 481706 14778 481942 15014
rect 481386 14458 481622 14694
rect 481706 14458 481942 14694
rect 481386 -3462 481622 -3226
rect 481706 -3462 481942 -3226
rect 481386 -3782 481622 -3546
rect 481706 -3782 481942 -3546
rect 485106 708442 485342 708678
rect 485426 708442 485662 708678
rect 485106 708122 485342 708358
rect 485426 708122 485662 708358
rect 485106 666498 485342 666734
rect 485426 666498 485662 666734
rect 485106 666178 485342 666414
rect 485426 666178 485662 666414
rect 485106 630498 485342 630734
rect 485426 630498 485662 630734
rect 485106 630178 485342 630414
rect 485426 630178 485662 630414
rect 485106 594498 485342 594734
rect 485426 594498 485662 594734
rect 485106 594178 485342 594414
rect 485426 594178 485662 594414
rect 485106 558498 485342 558734
rect 485426 558498 485662 558734
rect 485106 558178 485342 558414
rect 485426 558178 485662 558414
rect 485106 522498 485342 522734
rect 485426 522498 485662 522734
rect 485106 522178 485342 522414
rect 485426 522178 485662 522414
rect 485106 486498 485342 486734
rect 485426 486498 485662 486734
rect 485106 486178 485342 486414
rect 485426 486178 485662 486414
rect 485106 450498 485342 450734
rect 485426 450498 485662 450734
rect 485106 450178 485342 450414
rect 485426 450178 485662 450414
rect 485106 414498 485342 414734
rect 485426 414498 485662 414734
rect 485106 414178 485342 414414
rect 485426 414178 485662 414414
rect 485106 378498 485342 378734
rect 485426 378498 485662 378734
rect 485106 378178 485342 378414
rect 485426 378178 485662 378414
rect 485106 342498 485342 342734
rect 485426 342498 485662 342734
rect 485106 342178 485342 342414
rect 485426 342178 485662 342414
rect 485106 306498 485342 306734
rect 485426 306498 485662 306734
rect 485106 306178 485342 306414
rect 485426 306178 485662 306414
rect 485106 270498 485342 270734
rect 485426 270498 485662 270734
rect 485106 270178 485342 270414
rect 485426 270178 485662 270414
rect 485106 234498 485342 234734
rect 485426 234498 485662 234734
rect 485106 234178 485342 234414
rect 485426 234178 485662 234414
rect 485106 198498 485342 198734
rect 485426 198498 485662 198734
rect 485106 198178 485342 198414
rect 485426 198178 485662 198414
rect 485106 162498 485342 162734
rect 485426 162498 485662 162734
rect 485106 162178 485342 162414
rect 485426 162178 485662 162414
rect 485106 126498 485342 126734
rect 485426 126498 485662 126734
rect 485106 126178 485342 126414
rect 485426 126178 485662 126414
rect 485106 90498 485342 90734
rect 485426 90498 485662 90734
rect 485106 90178 485342 90414
rect 485426 90178 485662 90414
rect 485106 54498 485342 54734
rect 485426 54498 485662 54734
rect 485106 54178 485342 54414
rect 485426 54178 485662 54414
rect 485106 18498 485342 18734
rect 485426 18498 485662 18734
rect 485106 18178 485342 18414
rect 485426 18178 485662 18414
rect 485106 -4422 485342 -4186
rect 485426 -4422 485662 -4186
rect 485106 -4742 485342 -4506
rect 485426 -4742 485662 -4506
rect 488826 709402 489062 709638
rect 489146 709402 489382 709638
rect 488826 709082 489062 709318
rect 489146 709082 489382 709318
rect 488826 670218 489062 670454
rect 489146 670218 489382 670454
rect 488826 669898 489062 670134
rect 489146 669898 489382 670134
rect 488826 634218 489062 634454
rect 489146 634218 489382 634454
rect 488826 633898 489062 634134
rect 489146 633898 489382 634134
rect 488826 598218 489062 598454
rect 489146 598218 489382 598454
rect 488826 597898 489062 598134
rect 489146 597898 489382 598134
rect 488826 562218 489062 562454
rect 489146 562218 489382 562454
rect 488826 561898 489062 562134
rect 489146 561898 489382 562134
rect 488826 526218 489062 526454
rect 489146 526218 489382 526454
rect 488826 525898 489062 526134
rect 489146 525898 489382 526134
rect 488826 490218 489062 490454
rect 489146 490218 489382 490454
rect 488826 489898 489062 490134
rect 489146 489898 489382 490134
rect 488826 454218 489062 454454
rect 489146 454218 489382 454454
rect 488826 453898 489062 454134
rect 489146 453898 489382 454134
rect 488826 418218 489062 418454
rect 489146 418218 489382 418454
rect 488826 417898 489062 418134
rect 489146 417898 489382 418134
rect 488826 382218 489062 382454
rect 489146 382218 489382 382454
rect 488826 381898 489062 382134
rect 489146 381898 489382 382134
rect 488826 346218 489062 346454
rect 489146 346218 489382 346454
rect 488826 345898 489062 346134
rect 489146 345898 489382 346134
rect 488826 310218 489062 310454
rect 489146 310218 489382 310454
rect 488826 309898 489062 310134
rect 489146 309898 489382 310134
rect 488826 274218 489062 274454
rect 489146 274218 489382 274454
rect 488826 273898 489062 274134
rect 489146 273898 489382 274134
rect 488826 238218 489062 238454
rect 489146 238218 489382 238454
rect 488826 237898 489062 238134
rect 489146 237898 489382 238134
rect 488826 202218 489062 202454
rect 489146 202218 489382 202454
rect 488826 201898 489062 202134
rect 489146 201898 489382 202134
rect 488826 166218 489062 166454
rect 489146 166218 489382 166454
rect 488826 165898 489062 166134
rect 489146 165898 489382 166134
rect 488826 130218 489062 130454
rect 489146 130218 489382 130454
rect 488826 129898 489062 130134
rect 489146 129898 489382 130134
rect 488826 94218 489062 94454
rect 489146 94218 489382 94454
rect 488826 93898 489062 94134
rect 489146 93898 489382 94134
rect 488826 58218 489062 58454
rect 489146 58218 489382 58454
rect 488826 57898 489062 58134
rect 489146 57898 489382 58134
rect 488826 22218 489062 22454
rect 489146 22218 489382 22454
rect 488826 21898 489062 22134
rect 489146 21898 489382 22134
rect 488826 -5382 489062 -5146
rect 489146 -5382 489382 -5146
rect 488826 -5702 489062 -5466
rect 489146 -5702 489382 -5466
rect 492546 710362 492782 710598
rect 492866 710362 493102 710598
rect 492546 710042 492782 710278
rect 492866 710042 493102 710278
rect 492546 673938 492782 674174
rect 492866 673938 493102 674174
rect 492546 673618 492782 673854
rect 492866 673618 493102 673854
rect 492546 637938 492782 638174
rect 492866 637938 493102 638174
rect 492546 637618 492782 637854
rect 492866 637618 493102 637854
rect 492546 601938 492782 602174
rect 492866 601938 493102 602174
rect 492546 601618 492782 601854
rect 492866 601618 493102 601854
rect 492546 565938 492782 566174
rect 492866 565938 493102 566174
rect 492546 565618 492782 565854
rect 492866 565618 493102 565854
rect 492546 529938 492782 530174
rect 492866 529938 493102 530174
rect 492546 529618 492782 529854
rect 492866 529618 493102 529854
rect 492546 493938 492782 494174
rect 492866 493938 493102 494174
rect 492546 493618 492782 493854
rect 492866 493618 493102 493854
rect 492546 457938 492782 458174
rect 492866 457938 493102 458174
rect 492546 457618 492782 457854
rect 492866 457618 493102 457854
rect 492546 421938 492782 422174
rect 492866 421938 493102 422174
rect 492546 421618 492782 421854
rect 492866 421618 493102 421854
rect 492546 385938 492782 386174
rect 492866 385938 493102 386174
rect 492546 385618 492782 385854
rect 492866 385618 493102 385854
rect 492546 349938 492782 350174
rect 492866 349938 493102 350174
rect 492546 349618 492782 349854
rect 492866 349618 493102 349854
rect 492546 313938 492782 314174
rect 492866 313938 493102 314174
rect 492546 313618 492782 313854
rect 492866 313618 493102 313854
rect 492546 277938 492782 278174
rect 492866 277938 493102 278174
rect 492546 277618 492782 277854
rect 492866 277618 493102 277854
rect 492546 241938 492782 242174
rect 492866 241938 493102 242174
rect 492546 241618 492782 241854
rect 492866 241618 493102 241854
rect 492546 205938 492782 206174
rect 492866 205938 493102 206174
rect 492546 205618 492782 205854
rect 492866 205618 493102 205854
rect 492546 169938 492782 170174
rect 492866 169938 493102 170174
rect 492546 169618 492782 169854
rect 492866 169618 493102 169854
rect 492546 133938 492782 134174
rect 492866 133938 493102 134174
rect 492546 133618 492782 133854
rect 492866 133618 493102 133854
rect 492546 97938 492782 98174
rect 492866 97938 493102 98174
rect 492546 97618 492782 97854
rect 492866 97618 493102 97854
rect 492546 61938 492782 62174
rect 492866 61938 493102 62174
rect 492546 61618 492782 61854
rect 492866 61618 493102 61854
rect 492546 25938 492782 26174
rect 492866 25938 493102 26174
rect 492546 25618 492782 25854
rect 492866 25618 493102 25854
rect 492546 -6342 492782 -6106
rect 492866 -6342 493102 -6106
rect 492546 -6662 492782 -6426
rect 492866 -6662 493102 -6426
rect 496266 711322 496502 711558
rect 496586 711322 496822 711558
rect 496266 711002 496502 711238
rect 496586 711002 496822 711238
rect 496266 677658 496502 677894
rect 496586 677658 496822 677894
rect 496266 677338 496502 677574
rect 496586 677338 496822 677574
rect 496266 641658 496502 641894
rect 496586 641658 496822 641894
rect 496266 641338 496502 641574
rect 496586 641338 496822 641574
rect 496266 605658 496502 605894
rect 496586 605658 496822 605894
rect 496266 605338 496502 605574
rect 496586 605338 496822 605574
rect 496266 569658 496502 569894
rect 496586 569658 496822 569894
rect 496266 569338 496502 569574
rect 496586 569338 496822 569574
rect 496266 533658 496502 533894
rect 496586 533658 496822 533894
rect 496266 533338 496502 533574
rect 496586 533338 496822 533574
rect 496266 497658 496502 497894
rect 496586 497658 496822 497894
rect 496266 497338 496502 497574
rect 496586 497338 496822 497574
rect 496266 461658 496502 461894
rect 496586 461658 496822 461894
rect 496266 461338 496502 461574
rect 496586 461338 496822 461574
rect 496266 425658 496502 425894
rect 496586 425658 496822 425894
rect 496266 425338 496502 425574
rect 496586 425338 496822 425574
rect 496266 389658 496502 389894
rect 496586 389658 496822 389894
rect 496266 389338 496502 389574
rect 496586 389338 496822 389574
rect 496266 353658 496502 353894
rect 496586 353658 496822 353894
rect 496266 353338 496502 353574
rect 496586 353338 496822 353574
rect 496266 317658 496502 317894
rect 496586 317658 496822 317894
rect 496266 317338 496502 317574
rect 496586 317338 496822 317574
rect 496266 281658 496502 281894
rect 496586 281658 496822 281894
rect 496266 281338 496502 281574
rect 496586 281338 496822 281574
rect 496266 245658 496502 245894
rect 496586 245658 496822 245894
rect 496266 245338 496502 245574
rect 496586 245338 496822 245574
rect 496266 209658 496502 209894
rect 496586 209658 496822 209894
rect 496266 209338 496502 209574
rect 496586 209338 496822 209574
rect 496266 173658 496502 173894
rect 496586 173658 496822 173894
rect 496266 173338 496502 173574
rect 496586 173338 496822 173574
rect 496266 137658 496502 137894
rect 496586 137658 496822 137894
rect 496266 137338 496502 137574
rect 496586 137338 496822 137574
rect 496266 101658 496502 101894
rect 496586 101658 496822 101894
rect 496266 101338 496502 101574
rect 496586 101338 496822 101574
rect 496266 65658 496502 65894
rect 496586 65658 496822 65894
rect 496266 65338 496502 65574
rect 496586 65338 496822 65574
rect 496266 29658 496502 29894
rect 496586 29658 496822 29894
rect 496266 29338 496502 29574
rect 496586 29338 496822 29574
rect 496266 -7302 496502 -7066
rect 496586 -7302 496822 -7066
rect 496266 -7622 496502 -7386
rect 496586 -7622 496822 -7386
rect 506226 704602 506462 704838
rect 506546 704602 506782 704838
rect 506226 704282 506462 704518
rect 506546 704282 506782 704518
rect 506226 687618 506462 687854
rect 506546 687618 506782 687854
rect 506226 687298 506462 687534
rect 506546 687298 506782 687534
rect 506226 651618 506462 651854
rect 506546 651618 506782 651854
rect 506226 651298 506462 651534
rect 506546 651298 506782 651534
rect 506226 615618 506462 615854
rect 506546 615618 506782 615854
rect 506226 615298 506462 615534
rect 506546 615298 506782 615534
rect 506226 579618 506462 579854
rect 506546 579618 506782 579854
rect 506226 579298 506462 579534
rect 506546 579298 506782 579534
rect 506226 543618 506462 543854
rect 506546 543618 506782 543854
rect 506226 543298 506462 543534
rect 506546 543298 506782 543534
rect 506226 507618 506462 507854
rect 506546 507618 506782 507854
rect 506226 507298 506462 507534
rect 506546 507298 506782 507534
rect 506226 471618 506462 471854
rect 506546 471618 506782 471854
rect 506226 471298 506462 471534
rect 506546 471298 506782 471534
rect 506226 435618 506462 435854
rect 506546 435618 506782 435854
rect 506226 435298 506462 435534
rect 506546 435298 506782 435534
rect 506226 399618 506462 399854
rect 506546 399618 506782 399854
rect 506226 399298 506462 399534
rect 506546 399298 506782 399534
rect 506226 363618 506462 363854
rect 506546 363618 506782 363854
rect 506226 363298 506462 363534
rect 506546 363298 506782 363534
rect 506226 327618 506462 327854
rect 506546 327618 506782 327854
rect 506226 327298 506462 327534
rect 506546 327298 506782 327534
rect 506226 291618 506462 291854
rect 506546 291618 506782 291854
rect 506226 291298 506462 291534
rect 506546 291298 506782 291534
rect 506226 255618 506462 255854
rect 506546 255618 506782 255854
rect 506226 255298 506462 255534
rect 506546 255298 506782 255534
rect 506226 219618 506462 219854
rect 506546 219618 506782 219854
rect 506226 219298 506462 219534
rect 506546 219298 506782 219534
rect 506226 183618 506462 183854
rect 506546 183618 506782 183854
rect 506226 183298 506462 183534
rect 506546 183298 506782 183534
rect 506226 147618 506462 147854
rect 506546 147618 506782 147854
rect 506226 147298 506462 147534
rect 506546 147298 506782 147534
rect 506226 111618 506462 111854
rect 506546 111618 506782 111854
rect 506226 111298 506462 111534
rect 506546 111298 506782 111534
rect 506226 75618 506462 75854
rect 506546 75618 506782 75854
rect 506226 75298 506462 75534
rect 506546 75298 506782 75534
rect 506226 39618 506462 39854
rect 506546 39618 506782 39854
rect 506226 39298 506462 39534
rect 506546 39298 506782 39534
rect 506226 3618 506462 3854
rect 506546 3618 506782 3854
rect 506226 3298 506462 3534
rect 506546 3298 506782 3534
rect 506226 -582 506462 -346
rect 506546 -582 506782 -346
rect 506226 -902 506462 -666
rect 506546 -902 506782 -666
rect 509946 705562 510182 705798
rect 510266 705562 510502 705798
rect 509946 705242 510182 705478
rect 510266 705242 510502 705478
rect 509946 691338 510182 691574
rect 510266 691338 510502 691574
rect 509946 691018 510182 691254
rect 510266 691018 510502 691254
rect 509946 655338 510182 655574
rect 510266 655338 510502 655574
rect 509946 655018 510182 655254
rect 510266 655018 510502 655254
rect 509946 619338 510182 619574
rect 510266 619338 510502 619574
rect 509946 619018 510182 619254
rect 510266 619018 510502 619254
rect 509946 583338 510182 583574
rect 510266 583338 510502 583574
rect 509946 583018 510182 583254
rect 510266 583018 510502 583254
rect 509946 547338 510182 547574
rect 510266 547338 510502 547574
rect 509946 547018 510182 547254
rect 510266 547018 510502 547254
rect 509946 511338 510182 511574
rect 510266 511338 510502 511574
rect 509946 511018 510182 511254
rect 510266 511018 510502 511254
rect 509946 475338 510182 475574
rect 510266 475338 510502 475574
rect 509946 475018 510182 475254
rect 510266 475018 510502 475254
rect 509946 439338 510182 439574
rect 510266 439338 510502 439574
rect 509946 439018 510182 439254
rect 510266 439018 510502 439254
rect 509946 403338 510182 403574
rect 510266 403338 510502 403574
rect 509946 403018 510182 403254
rect 510266 403018 510502 403254
rect 509946 367338 510182 367574
rect 510266 367338 510502 367574
rect 509946 367018 510182 367254
rect 510266 367018 510502 367254
rect 509946 331338 510182 331574
rect 510266 331338 510502 331574
rect 509946 331018 510182 331254
rect 510266 331018 510502 331254
rect 509946 295338 510182 295574
rect 510266 295338 510502 295574
rect 509946 295018 510182 295254
rect 510266 295018 510502 295254
rect 509946 259338 510182 259574
rect 510266 259338 510502 259574
rect 509946 259018 510182 259254
rect 510266 259018 510502 259254
rect 509946 223338 510182 223574
rect 510266 223338 510502 223574
rect 509946 223018 510182 223254
rect 510266 223018 510502 223254
rect 509946 187338 510182 187574
rect 510266 187338 510502 187574
rect 509946 187018 510182 187254
rect 510266 187018 510502 187254
rect 509946 151338 510182 151574
rect 510266 151338 510502 151574
rect 509946 151018 510182 151254
rect 510266 151018 510502 151254
rect 509946 115338 510182 115574
rect 510266 115338 510502 115574
rect 509946 115018 510182 115254
rect 510266 115018 510502 115254
rect 509946 79338 510182 79574
rect 510266 79338 510502 79574
rect 509946 79018 510182 79254
rect 510266 79018 510502 79254
rect 509946 43338 510182 43574
rect 510266 43338 510502 43574
rect 509946 43018 510182 43254
rect 510266 43018 510502 43254
rect 509946 7338 510182 7574
rect 510266 7338 510502 7574
rect 509946 7018 510182 7254
rect 510266 7018 510502 7254
rect 509946 -1542 510182 -1306
rect 510266 -1542 510502 -1306
rect 509946 -1862 510182 -1626
rect 510266 -1862 510502 -1626
rect 513666 706522 513902 706758
rect 513986 706522 514222 706758
rect 513666 706202 513902 706438
rect 513986 706202 514222 706438
rect 513666 695058 513902 695294
rect 513986 695058 514222 695294
rect 513666 694738 513902 694974
rect 513986 694738 514222 694974
rect 513666 659058 513902 659294
rect 513986 659058 514222 659294
rect 513666 658738 513902 658974
rect 513986 658738 514222 658974
rect 513666 623058 513902 623294
rect 513986 623058 514222 623294
rect 513666 622738 513902 622974
rect 513986 622738 514222 622974
rect 513666 587058 513902 587294
rect 513986 587058 514222 587294
rect 513666 586738 513902 586974
rect 513986 586738 514222 586974
rect 513666 551058 513902 551294
rect 513986 551058 514222 551294
rect 513666 550738 513902 550974
rect 513986 550738 514222 550974
rect 513666 515058 513902 515294
rect 513986 515058 514222 515294
rect 513666 514738 513902 514974
rect 513986 514738 514222 514974
rect 513666 479058 513902 479294
rect 513986 479058 514222 479294
rect 513666 478738 513902 478974
rect 513986 478738 514222 478974
rect 513666 443058 513902 443294
rect 513986 443058 514222 443294
rect 513666 442738 513902 442974
rect 513986 442738 514222 442974
rect 513666 407058 513902 407294
rect 513986 407058 514222 407294
rect 513666 406738 513902 406974
rect 513986 406738 514222 406974
rect 513666 371058 513902 371294
rect 513986 371058 514222 371294
rect 513666 370738 513902 370974
rect 513986 370738 514222 370974
rect 513666 335058 513902 335294
rect 513986 335058 514222 335294
rect 513666 334738 513902 334974
rect 513986 334738 514222 334974
rect 513666 299058 513902 299294
rect 513986 299058 514222 299294
rect 513666 298738 513902 298974
rect 513986 298738 514222 298974
rect 513666 263058 513902 263294
rect 513986 263058 514222 263294
rect 513666 262738 513902 262974
rect 513986 262738 514222 262974
rect 513666 227058 513902 227294
rect 513986 227058 514222 227294
rect 513666 226738 513902 226974
rect 513986 226738 514222 226974
rect 513666 191058 513902 191294
rect 513986 191058 514222 191294
rect 513666 190738 513902 190974
rect 513986 190738 514222 190974
rect 513666 155058 513902 155294
rect 513986 155058 514222 155294
rect 513666 154738 513902 154974
rect 513986 154738 514222 154974
rect 513666 119058 513902 119294
rect 513986 119058 514222 119294
rect 513666 118738 513902 118974
rect 513986 118738 514222 118974
rect 513666 83058 513902 83294
rect 513986 83058 514222 83294
rect 513666 82738 513902 82974
rect 513986 82738 514222 82974
rect 513666 47058 513902 47294
rect 513986 47058 514222 47294
rect 513666 46738 513902 46974
rect 513986 46738 514222 46974
rect 513666 11058 513902 11294
rect 513986 11058 514222 11294
rect 513666 10738 513902 10974
rect 513986 10738 514222 10974
rect 513666 -2502 513902 -2266
rect 513986 -2502 514222 -2266
rect 513666 -2822 513902 -2586
rect 513986 -2822 514222 -2586
rect 517386 707482 517622 707718
rect 517706 707482 517942 707718
rect 517386 707162 517622 707398
rect 517706 707162 517942 707398
rect 517386 698778 517622 699014
rect 517706 698778 517942 699014
rect 517386 698458 517622 698694
rect 517706 698458 517942 698694
rect 517386 662778 517622 663014
rect 517706 662778 517942 663014
rect 517386 662458 517622 662694
rect 517706 662458 517942 662694
rect 517386 626778 517622 627014
rect 517706 626778 517942 627014
rect 517386 626458 517622 626694
rect 517706 626458 517942 626694
rect 517386 590778 517622 591014
rect 517706 590778 517942 591014
rect 517386 590458 517622 590694
rect 517706 590458 517942 590694
rect 517386 554778 517622 555014
rect 517706 554778 517942 555014
rect 517386 554458 517622 554694
rect 517706 554458 517942 554694
rect 517386 518778 517622 519014
rect 517706 518778 517942 519014
rect 517386 518458 517622 518694
rect 517706 518458 517942 518694
rect 517386 482778 517622 483014
rect 517706 482778 517942 483014
rect 517386 482458 517622 482694
rect 517706 482458 517942 482694
rect 517386 446778 517622 447014
rect 517706 446778 517942 447014
rect 517386 446458 517622 446694
rect 517706 446458 517942 446694
rect 517386 410778 517622 411014
rect 517706 410778 517942 411014
rect 517386 410458 517622 410694
rect 517706 410458 517942 410694
rect 517386 374778 517622 375014
rect 517706 374778 517942 375014
rect 517386 374458 517622 374694
rect 517706 374458 517942 374694
rect 517386 338778 517622 339014
rect 517706 338778 517942 339014
rect 517386 338458 517622 338694
rect 517706 338458 517942 338694
rect 517386 302778 517622 303014
rect 517706 302778 517942 303014
rect 517386 302458 517622 302694
rect 517706 302458 517942 302694
rect 517386 266778 517622 267014
rect 517706 266778 517942 267014
rect 517386 266458 517622 266694
rect 517706 266458 517942 266694
rect 517386 230778 517622 231014
rect 517706 230778 517942 231014
rect 517386 230458 517622 230694
rect 517706 230458 517942 230694
rect 517386 194778 517622 195014
rect 517706 194778 517942 195014
rect 517386 194458 517622 194694
rect 517706 194458 517942 194694
rect 517386 158778 517622 159014
rect 517706 158778 517942 159014
rect 517386 158458 517622 158694
rect 517706 158458 517942 158694
rect 517386 122778 517622 123014
rect 517706 122778 517942 123014
rect 517386 122458 517622 122694
rect 517706 122458 517942 122694
rect 517386 86778 517622 87014
rect 517706 86778 517942 87014
rect 517386 86458 517622 86694
rect 517706 86458 517942 86694
rect 517386 50778 517622 51014
rect 517706 50778 517942 51014
rect 517386 50458 517622 50694
rect 517706 50458 517942 50694
rect 517386 14778 517622 15014
rect 517706 14778 517942 15014
rect 517386 14458 517622 14694
rect 517706 14458 517942 14694
rect 517386 -3462 517622 -3226
rect 517706 -3462 517942 -3226
rect 517386 -3782 517622 -3546
rect 517706 -3782 517942 -3546
rect 521106 708442 521342 708678
rect 521426 708442 521662 708678
rect 521106 708122 521342 708358
rect 521426 708122 521662 708358
rect 521106 666498 521342 666734
rect 521426 666498 521662 666734
rect 521106 666178 521342 666414
rect 521426 666178 521662 666414
rect 521106 630498 521342 630734
rect 521426 630498 521662 630734
rect 521106 630178 521342 630414
rect 521426 630178 521662 630414
rect 521106 594498 521342 594734
rect 521426 594498 521662 594734
rect 521106 594178 521342 594414
rect 521426 594178 521662 594414
rect 521106 558498 521342 558734
rect 521426 558498 521662 558734
rect 521106 558178 521342 558414
rect 521426 558178 521662 558414
rect 521106 522498 521342 522734
rect 521426 522498 521662 522734
rect 521106 522178 521342 522414
rect 521426 522178 521662 522414
rect 521106 486498 521342 486734
rect 521426 486498 521662 486734
rect 521106 486178 521342 486414
rect 521426 486178 521662 486414
rect 521106 450498 521342 450734
rect 521426 450498 521662 450734
rect 521106 450178 521342 450414
rect 521426 450178 521662 450414
rect 521106 414498 521342 414734
rect 521426 414498 521662 414734
rect 521106 414178 521342 414414
rect 521426 414178 521662 414414
rect 521106 378498 521342 378734
rect 521426 378498 521662 378734
rect 521106 378178 521342 378414
rect 521426 378178 521662 378414
rect 521106 342498 521342 342734
rect 521426 342498 521662 342734
rect 521106 342178 521342 342414
rect 521426 342178 521662 342414
rect 521106 306498 521342 306734
rect 521426 306498 521662 306734
rect 521106 306178 521342 306414
rect 521426 306178 521662 306414
rect 521106 270498 521342 270734
rect 521426 270498 521662 270734
rect 521106 270178 521342 270414
rect 521426 270178 521662 270414
rect 521106 234498 521342 234734
rect 521426 234498 521662 234734
rect 521106 234178 521342 234414
rect 521426 234178 521662 234414
rect 521106 198498 521342 198734
rect 521426 198498 521662 198734
rect 521106 198178 521342 198414
rect 521426 198178 521662 198414
rect 521106 162498 521342 162734
rect 521426 162498 521662 162734
rect 521106 162178 521342 162414
rect 521426 162178 521662 162414
rect 521106 126498 521342 126734
rect 521426 126498 521662 126734
rect 521106 126178 521342 126414
rect 521426 126178 521662 126414
rect 521106 90498 521342 90734
rect 521426 90498 521662 90734
rect 521106 90178 521342 90414
rect 521426 90178 521662 90414
rect 521106 54498 521342 54734
rect 521426 54498 521662 54734
rect 521106 54178 521342 54414
rect 521426 54178 521662 54414
rect 521106 18498 521342 18734
rect 521426 18498 521662 18734
rect 521106 18178 521342 18414
rect 521426 18178 521662 18414
rect 521106 -4422 521342 -4186
rect 521426 -4422 521662 -4186
rect 521106 -4742 521342 -4506
rect 521426 -4742 521662 -4506
rect 524826 709402 525062 709638
rect 525146 709402 525382 709638
rect 524826 709082 525062 709318
rect 525146 709082 525382 709318
rect 524826 670218 525062 670454
rect 525146 670218 525382 670454
rect 524826 669898 525062 670134
rect 525146 669898 525382 670134
rect 524826 634218 525062 634454
rect 525146 634218 525382 634454
rect 524826 633898 525062 634134
rect 525146 633898 525382 634134
rect 524826 598218 525062 598454
rect 525146 598218 525382 598454
rect 524826 597898 525062 598134
rect 525146 597898 525382 598134
rect 524826 562218 525062 562454
rect 525146 562218 525382 562454
rect 524826 561898 525062 562134
rect 525146 561898 525382 562134
rect 524826 526218 525062 526454
rect 525146 526218 525382 526454
rect 524826 525898 525062 526134
rect 525146 525898 525382 526134
rect 524826 490218 525062 490454
rect 525146 490218 525382 490454
rect 524826 489898 525062 490134
rect 525146 489898 525382 490134
rect 524826 454218 525062 454454
rect 525146 454218 525382 454454
rect 524826 453898 525062 454134
rect 525146 453898 525382 454134
rect 524826 418218 525062 418454
rect 525146 418218 525382 418454
rect 524826 417898 525062 418134
rect 525146 417898 525382 418134
rect 524826 382218 525062 382454
rect 525146 382218 525382 382454
rect 524826 381898 525062 382134
rect 525146 381898 525382 382134
rect 524826 346218 525062 346454
rect 525146 346218 525382 346454
rect 524826 345898 525062 346134
rect 525146 345898 525382 346134
rect 524826 310218 525062 310454
rect 525146 310218 525382 310454
rect 524826 309898 525062 310134
rect 525146 309898 525382 310134
rect 524826 274218 525062 274454
rect 525146 274218 525382 274454
rect 524826 273898 525062 274134
rect 525146 273898 525382 274134
rect 524826 238218 525062 238454
rect 525146 238218 525382 238454
rect 524826 237898 525062 238134
rect 525146 237898 525382 238134
rect 524826 202218 525062 202454
rect 525146 202218 525382 202454
rect 524826 201898 525062 202134
rect 525146 201898 525382 202134
rect 524826 166218 525062 166454
rect 525146 166218 525382 166454
rect 524826 165898 525062 166134
rect 525146 165898 525382 166134
rect 524826 130218 525062 130454
rect 525146 130218 525382 130454
rect 524826 129898 525062 130134
rect 525146 129898 525382 130134
rect 524826 94218 525062 94454
rect 525146 94218 525382 94454
rect 524826 93898 525062 94134
rect 525146 93898 525382 94134
rect 524826 58218 525062 58454
rect 525146 58218 525382 58454
rect 524826 57898 525062 58134
rect 525146 57898 525382 58134
rect 524826 22218 525062 22454
rect 525146 22218 525382 22454
rect 524826 21898 525062 22134
rect 525146 21898 525382 22134
rect 524826 -5382 525062 -5146
rect 525146 -5382 525382 -5146
rect 524826 -5702 525062 -5466
rect 525146 -5702 525382 -5466
rect 528546 710362 528782 710598
rect 528866 710362 529102 710598
rect 528546 710042 528782 710278
rect 528866 710042 529102 710278
rect 528546 673938 528782 674174
rect 528866 673938 529102 674174
rect 528546 673618 528782 673854
rect 528866 673618 529102 673854
rect 528546 637938 528782 638174
rect 528866 637938 529102 638174
rect 528546 637618 528782 637854
rect 528866 637618 529102 637854
rect 528546 601938 528782 602174
rect 528866 601938 529102 602174
rect 528546 601618 528782 601854
rect 528866 601618 529102 601854
rect 528546 565938 528782 566174
rect 528866 565938 529102 566174
rect 528546 565618 528782 565854
rect 528866 565618 529102 565854
rect 528546 529938 528782 530174
rect 528866 529938 529102 530174
rect 528546 529618 528782 529854
rect 528866 529618 529102 529854
rect 528546 493938 528782 494174
rect 528866 493938 529102 494174
rect 528546 493618 528782 493854
rect 528866 493618 529102 493854
rect 528546 457938 528782 458174
rect 528866 457938 529102 458174
rect 528546 457618 528782 457854
rect 528866 457618 529102 457854
rect 528546 421938 528782 422174
rect 528866 421938 529102 422174
rect 528546 421618 528782 421854
rect 528866 421618 529102 421854
rect 528546 385938 528782 386174
rect 528866 385938 529102 386174
rect 528546 385618 528782 385854
rect 528866 385618 529102 385854
rect 528546 349938 528782 350174
rect 528866 349938 529102 350174
rect 528546 349618 528782 349854
rect 528866 349618 529102 349854
rect 528546 313938 528782 314174
rect 528866 313938 529102 314174
rect 528546 313618 528782 313854
rect 528866 313618 529102 313854
rect 528546 277938 528782 278174
rect 528866 277938 529102 278174
rect 528546 277618 528782 277854
rect 528866 277618 529102 277854
rect 528546 241938 528782 242174
rect 528866 241938 529102 242174
rect 528546 241618 528782 241854
rect 528866 241618 529102 241854
rect 528546 205938 528782 206174
rect 528866 205938 529102 206174
rect 528546 205618 528782 205854
rect 528866 205618 529102 205854
rect 528546 169938 528782 170174
rect 528866 169938 529102 170174
rect 528546 169618 528782 169854
rect 528866 169618 529102 169854
rect 528546 133938 528782 134174
rect 528866 133938 529102 134174
rect 528546 133618 528782 133854
rect 528866 133618 529102 133854
rect 528546 97938 528782 98174
rect 528866 97938 529102 98174
rect 528546 97618 528782 97854
rect 528866 97618 529102 97854
rect 528546 61938 528782 62174
rect 528866 61938 529102 62174
rect 528546 61618 528782 61854
rect 528866 61618 529102 61854
rect 528546 25938 528782 26174
rect 528866 25938 529102 26174
rect 528546 25618 528782 25854
rect 528866 25618 529102 25854
rect 528546 -6342 528782 -6106
rect 528866 -6342 529102 -6106
rect 528546 -6662 528782 -6426
rect 528866 -6662 529102 -6426
rect 532266 711322 532502 711558
rect 532586 711322 532822 711558
rect 532266 711002 532502 711238
rect 532586 711002 532822 711238
rect 532266 677658 532502 677894
rect 532586 677658 532822 677894
rect 532266 677338 532502 677574
rect 532586 677338 532822 677574
rect 532266 641658 532502 641894
rect 532586 641658 532822 641894
rect 532266 641338 532502 641574
rect 532586 641338 532822 641574
rect 532266 605658 532502 605894
rect 532586 605658 532822 605894
rect 532266 605338 532502 605574
rect 532586 605338 532822 605574
rect 532266 569658 532502 569894
rect 532586 569658 532822 569894
rect 532266 569338 532502 569574
rect 532586 569338 532822 569574
rect 532266 533658 532502 533894
rect 532586 533658 532822 533894
rect 532266 533338 532502 533574
rect 532586 533338 532822 533574
rect 532266 497658 532502 497894
rect 532586 497658 532822 497894
rect 532266 497338 532502 497574
rect 532586 497338 532822 497574
rect 532266 461658 532502 461894
rect 532586 461658 532822 461894
rect 532266 461338 532502 461574
rect 532586 461338 532822 461574
rect 532266 425658 532502 425894
rect 532586 425658 532822 425894
rect 532266 425338 532502 425574
rect 532586 425338 532822 425574
rect 532266 389658 532502 389894
rect 532586 389658 532822 389894
rect 532266 389338 532502 389574
rect 532586 389338 532822 389574
rect 532266 353658 532502 353894
rect 532586 353658 532822 353894
rect 532266 353338 532502 353574
rect 532586 353338 532822 353574
rect 532266 317658 532502 317894
rect 532586 317658 532822 317894
rect 532266 317338 532502 317574
rect 532586 317338 532822 317574
rect 532266 281658 532502 281894
rect 532586 281658 532822 281894
rect 532266 281338 532502 281574
rect 532586 281338 532822 281574
rect 532266 245658 532502 245894
rect 532586 245658 532822 245894
rect 532266 245338 532502 245574
rect 532586 245338 532822 245574
rect 532266 209658 532502 209894
rect 532586 209658 532822 209894
rect 532266 209338 532502 209574
rect 532586 209338 532822 209574
rect 532266 173658 532502 173894
rect 532586 173658 532822 173894
rect 532266 173338 532502 173574
rect 532586 173338 532822 173574
rect 532266 137658 532502 137894
rect 532586 137658 532822 137894
rect 532266 137338 532502 137574
rect 532586 137338 532822 137574
rect 532266 101658 532502 101894
rect 532586 101658 532822 101894
rect 532266 101338 532502 101574
rect 532586 101338 532822 101574
rect 532266 65658 532502 65894
rect 532586 65658 532822 65894
rect 532266 65338 532502 65574
rect 532586 65338 532822 65574
rect 532266 29658 532502 29894
rect 532586 29658 532822 29894
rect 532266 29338 532502 29574
rect 532586 29338 532822 29574
rect 532266 -7302 532502 -7066
rect 532586 -7302 532822 -7066
rect 532266 -7622 532502 -7386
rect 532586 -7622 532822 -7386
rect 542226 704602 542462 704838
rect 542546 704602 542782 704838
rect 542226 704282 542462 704518
rect 542546 704282 542782 704518
rect 542226 687618 542462 687854
rect 542546 687618 542782 687854
rect 542226 687298 542462 687534
rect 542546 687298 542782 687534
rect 542226 651618 542462 651854
rect 542546 651618 542782 651854
rect 542226 651298 542462 651534
rect 542546 651298 542782 651534
rect 542226 615618 542462 615854
rect 542546 615618 542782 615854
rect 542226 615298 542462 615534
rect 542546 615298 542782 615534
rect 542226 579618 542462 579854
rect 542546 579618 542782 579854
rect 542226 579298 542462 579534
rect 542546 579298 542782 579534
rect 542226 543618 542462 543854
rect 542546 543618 542782 543854
rect 542226 543298 542462 543534
rect 542546 543298 542782 543534
rect 542226 507618 542462 507854
rect 542546 507618 542782 507854
rect 542226 507298 542462 507534
rect 542546 507298 542782 507534
rect 542226 471618 542462 471854
rect 542546 471618 542782 471854
rect 542226 471298 542462 471534
rect 542546 471298 542782 471534
rect 542226 435618 542462 435854
rect 542546 435618 542782 435854
rect 542226 435298 542462 435534
rect 542546 435298 542782 435534
rect 542226 399618 542462 399854
rect 542546 399618 542782 399854
rect 542226 399298 542462 399534
rect 542546 399298 542782 399534
rect 542226 363618 542462 363854
rect 542546 363618 542782 363854
rect 542226 363298 542462 363534
rect 542546 363298 542782 363534
rect 542226 327618 542462 327854
rect 542546 327618 542782 327854
rect 542226 327298 542462 327534
rect 542546 327298 542782 327534
rect 542226 291618 542462 291854
rect 542546 291618 542782 291854
rect 542226 291298 542462 291534
rect 542546 291298 542782 291534
rect 542226 255618 542462 255854
rect 542546 255618 542782 255854
rect 542226 255298 542462 255534
rect 542546 255298 542782 255534
rect 542226 219618 542462 219854
rect 542546 219618 542782 219854
rect 542226 219298 542462 219534
rect 542546 219298 542782 219534
rect 542226 183618 542462 183854
rect 542546 183618 542782 183854
rect 542226 183298 542462 183534
rect 542546 183298 542782 183534
rect 542226 147618 542462 147854
rect 542546 147618 542782 147854
rect 542226 147298 542462 147534
rect 542546 147298 542782 147534
rect 542226 111618 542462 111854
rect 542546 111618 542782 111854
rect 542226 111298 542462 111534
rect 542546 111298 542782 111534
rect 542226 75618 542462 75854
rect 542546 75618 542782 75854
rect 542226 75298 542462 75534
rect 542546 75298 542782 75534
rect 542226 39618 542462 39854
rect 542546 39618 542782 39854
rect 542226 39298 542462 39534
rect 542546 39298 542782 39534
rect 542226 3618 542462 3854
rect 542546 3618 542782 3854
rect 542226 3298 542462 3534
rect 542546 3298 542782 3534
rect 542226 -582 542462 -346
rect 542546 -582 542782 -346
rect 542226 -902 542462 -666
rect 542546 -902 542782 -666
rect 545946 705562 546182 705798
rect 546266 705562 546502 705798
rect 545946 705242 546182 705478
rect 546266 705242 546502 705478
rect 545946 691338 546182 691574
rect 546266 691338 546502 691574
rect 545946 691018 546182 691254
rect 546266 691018 546502 691254
rect 545946 655338 546182 655574
rect 546266 655338 546502 655574
rect 545946 655018 546182 655254
rect 546266 655018 546502 655254
rect 545946 619338 546182 619574
rect 546266 619338 546502 619574
rect 545946 619018 546182 619254
rect 546266 619018 546502 619254
rect 545946 583338 546182 583574
rect 546266 583338 546502 583574
rect 545946 583018 546182 583254
rect 546266 583018 546502 583254
rect 545946 547338 546182 547574
rect 546266 547338 546502 547574
rect 545946 547018 546182 547254
rect 546266 547018 546502 547254
rect 545946 511338 546182 511574
rect 546266 511338 546502 511574
rect 545946 511018 546182 511254
rect 546266 511018 546502 511254
rect 545946 475338 546182 475574
rect 546266 475338 546502 475574
rect 545946 475018 546182 475254
rect 546266 475018 546502 475254
rect 545946 439338 546182 439574
rect 546266 439338 546502 439574
rect 545946 439018 546182 439254
rect 546266 439018 546502 439254
rect 545946 403338 546182 403574
rect 546266 403338 546502 403574
rect 545946 403018 546182 403254
rect 546266 403018 546502 403254
rect 545946 367338 546182 367574
rect 546266 367338 546502 367574
rect 545946 367018 546182 367254
rect 546266 367018 546502 367254
rect 545946 331338 546182 331574
rect 546266 331338 546502 331574
rect 545946 331018 546182 331254
rect 546266 331018 546502 331254
rect 545946 295338 546182 295574
rect 546266 295338 546502 295574
rect 545946 295018 546182 295254
rect 546266 295018 546502 295254
rect 545946 259338 546182 259574
rect 546266 259338 546502 259574
rect 545946 259018 546182 259254
rect 546266 259018 546502 259254
rect 545946 223338 546182 223574
rect 546266 223338 546502 223574
rect 545946 223018 546182 223254
rect 546266 223018 546502 223254
rect 545946 187338 546182 187574
rect 546266 187338 546502 187574
rect 545946 187018 546182 187254
rect 546266 187018 546502 187254
rect 545946 151338 546182 151574
rect 546266 151338 546502 151574
rect 545946 151018 546182 151254
rect 546266 151018 546502 151254
rect 545946 115338 546182 115574
rect 546266 115338 546502 115574
rect 545946 115018 546182 115254
rect 546266 115018 546502 115254
rect 545946 79338 546182 79574
rect 546266 79338 546502 79574
rect 545946 79018 546182 79254
rect 546266 79018 546502 79254
rect 545946 43338 546182 43574
rect 546266 43338 546502 43574
rect 545946 43018 546182 43254
rect 546266 43018 546502 43254
rect 545946 7338 546182 7574
rect 546266 7338 546502 7574
rect 545946 7018 546182 7254
rect 546266 7018 546502 7254
rect 545946 -1542 546182 -1306
rect 546266 -1542 546502 -1306
rect 545946 -1862 546182 -1626
rect 546266 -1862 546502 -1626
rect 549666 706522 549902 706758
rect 549986 706522 550222 706758
rect 549666 706202 549902 706438
rect 549986 706202 550222 706438
rect 549666 695058 549902 695294
rect 549986 695058 550222 695294
rect 549666 694738 549902 694974
rect 549986 694738 550222 694974
rect 549666 659058 549902 659294
rect 549986 659058 550222 659294
rect 549666 658738 549902 658974
rect 549986 658738 550222 658974
rect 549666 623058 549902 623294
rect 549986 623058 550222 623294
rect 549666 622738 549902 622974
rect 549986 622738 550222 622974
rect 549666 587058 549902 587294
rect 549986 587058 550222 587294
rect 549666 586738 549902 586974
rect 549986 586738 550222 586974
rect 549666 551058 549902 551294
rect 549986 551058 550222 551294
rect 549666 550738 549902 550974
rect 549986 550738 550222 550974
rect 549666 515058 549902 515294
rect 549986 515058 550222 515294
rect 549666 514738 549902 514974
rect 549986 514738 550222 514974
rect 549666 479058 549902 479294
rect 549986 479058 550222 479294
rect 549666 478738 549902 478974
rect 549986 478738 550222 478974
rect 549666 443058 549902 443294
rect 549986 443058 550222 443294
rect 549666 442738 549902 442974
rect 549986 442738 550222 442974
rect 549666 407058 549902 407294
rect 549986 407058 550222 407294
rect 549666 406738 549902 406974
rect 549986 406738 550222 406974
rect 549666 371058 549902 371294
rect 549986 371058 550222 371294
rect 549666 370738 549902 370974
rect 549986 370738 550222 370974
rect 549666 335058 549902 335294
rect 549986 335058 550222 335294
rect 549666 334738 549902 334974
rect 549986 334738 550222 334974
rect 549666 299058 549902 299294
rect 549986 299058 550222 299294
rect 549666 298738 549902 298974
rect 549986 298738 550222 298974
rect 549666 263058 549902 263294
rect 549986 263058 550222 263294
rect 549666 262738 549902 262974
rect 549986 262738 550222 262974
rect 549666 227058 549902 227294
rect 549986 227058 550222 227294
rect 549666 226738 549902 226974
rect 549986 226738 550222 226974
rect 549666 191058 549902 191294
rect 549986 191058 550222 191294
rect 549666 190738 549902 190974
rect 549986 190738 550222 190974
rect 549666 155058 549902 155294
rect 549986 155058 550222 155294
rect 549666 154738 549902 154974
rect 549986 154738 550222 154974
rect 549666 119058 549902 119294
rect 549986 119058 550222 119294
rect 549666 118738 549902 118974
rect 549986 118738 550222 118974
rect 549666 83058 549902 83294
rect 549986 83058 550222 83294
rect 549666 82738 549902 82974
rect 549986 82738 550222 82974
rect 549666 47058 549902 47294
rect 549986 47058 550222 47294
rect 549666 46738 549902 46974
rect 549986 46738 550222 46974
rect 549666 11058 549902 11294
rect 549986 11058 550222 11294
rect 549666 10738 549902 10974
rect 549986 10738 550222 10974
rect 549666 -2502 549902 -2266
rect 549986 -2502 550222 -2266
rect 549666 -2822 549902 -2586
rect 549986 -2822 550222 -2586
rect 553386 707482 553622 707718
rect 553706 707482 553942 707718
rect 553386 707162 553622 707398
rect 553706 707162 553942 707398
rect 553386 698778 553622 699014
rect 553706 698778 553942 699014
rect 553386 698458 553622 698694
rect 553706 698458 553942 698694
rect 553386 662778 553622 663014
rect 553706 662778 553942 663014
rect 553386 662458 553622 662694
rect 553706 662458 553942 662694
rect 553386 626778 553622 627014
rect 553706 626778 553942 627014
rect 553386 626458 553622 626694
rect 553706 626458 553942 626694
rect 553386 590778 553622 591014
rect 553706 590778 553942 591014
rect 553386 590458 553622 590694
rect 553706 590458 553942 590694
rect 553386 554778 553622 555014
rect 553706 554778 553942 555014
rect 553386 554458 553622 554694
rect 553706 554458 553942 554694
rect 553386 518778 553622 519014
rect 553706 518778 553942 519014
rect 553386 518458 553622 518694
rect 553706 518458 553942 518694
rect 553386 482778 553622 483014
rect 553706 482778 553942 483014
rect 553386 482458 553622 482694
rect 553706 482458 553942 482694
rect 553386 446778 553622 447014
rect 553706 446778 553942 447014
rect 553386 446458 553622 446694
rect 553706 446458 553942 446694
rect 553386 410778 553622 411014
rect 553706 410778 553942 411014
rect 553386 410458 553622 410694
rect 553706 410458 553942 410694
rect 553386 374778 553622 375014
rect 553706 374778 553942 375014
rect 553386 374458 553622 374694
rect 553706 374458 553942 374694
rect 553386 338778 553622 339014
rect 553706 338778 553942 339014
rect 553386 338458 553622 338694
rect 553706 338458 553942 338694
rect 553386 302778 553622 303014
rect 553706 302778 553942 303014
rect 553386 302458 553622 302694
rect 553706 302458 553942 302694
rect 553386 266778 553622 267014
rect 553706 266778 553942 267014
rect 553386 266458 553622 266694
rect 553706 266458 553942 266694
rect 553386 230778 553622 231014
rect 553706 230778 553942 231014
rect 553386 230458 553622 230694
rect 553706 230458 553942 230694
rect 553386 194778 553622 195014
rect 553706 194778 553942 195014
rect 553386 194458 553622 194694
rect 553706 194458 553942 194694
rect 553386 158778 553622 159014
rect 553706 158778 553942 159014
rect 553386 158458 553622 158694
rect 553706 158458 553942 158694
rect 553386 122778 553622 123014
rect 553706 122778 553942 123014
rect 553386 122458 553622 122694
rect 553706 122458 553942 122694
rect 553386 86778 553622 87014
rect 553706 86778 553942 87014
rect 553386 86458 553622 86694
rect 553706 86458 553942 86694
rect 553386 50778 553622 51014
rect 553706 50778 553942 51014
rect 553386 50458 553622 50694
rect 553706 50458 553942 50694
rect 553386 14778 553622 15014
rect 553706 14778 553942 15014
rect 553386 14458 553622 14694
rect 553706 14458 553942 14694
rect 553386 -3462 553622 -3226
rect 553706 -3462 553942 -3226
rect 553386 -3782 553622 -3546
rect 553706 -3782 553942 -3546
rect 557106 708442 557342 708678
rect 557426 708442 557662 708678
rect 557106 708122 557342 708358
rect 557426 708122 557662 708358
rect 557106 666498 557342 666734
rect 557426 666498 557662 666734
rect 557106 666178 557342 666414
rect 557426 666178 557662 666414
rect 557106 630498 557342 630734
rect 557426 630498 557662 630734
rect 557106 630178 557342 630414
rect 557426 630178 557662 630414
rect 557106 594498 557342 594734
rect 557426 594498 557662 594734
rect 557106 594178 557342 594414
rect 557426 594178 557662 594414
rect 557106 558498 557342 558734
rect 557426 558498 557662 558734
rect 557106 558178 557342 558414
rect 557426 558178 557662 558414
rect 557106 522498 557342 522734
rect 557426 522498 557662 522734
rect 557106 522178 557342 522414
rect 557426 522178 557662 522414
rect 557106 486498 557342 486734
rect 557426 486498 557662 486734
rect 557106 486178 557342 486414
rect 557426 486178 557662 486414
rect 557106 450498 557342 450734
rect 557426 450498 557662 450734
rect 557106 450178 557342 450414
rect 557426 450178 557662 450414
rect 557106 414498 557342 414734
rect 557426 414498 557662 414734
rect 557106 414178 557342 414414
rect 557426 414178 557662 414414
rect 557106 378498 557342 378734
rect 557426 378498 557662 378734
rect 557106 378178 557342 378414
rect 557426 378178 557662 378414
rect 557106 342498 557342 342734
rect 557426 342498 557662 342734
rect 557106 342178 557342 342414
rect 557426 342178 557662 342414
rect 557106 306498 557342 306734
rect 557426 306498 557662 306734
rect 557106 306178 557342 306414
rect 557426 306178 557662 306414
rect 557106 270498 557342 270734
rect 557426 270498 557662 270734
rect 557106 270178 557342 270414
rect 557426 270178 557662 270414
rect 557106 234498 557342 234734
rect 557426 234498 557662 234734
rect 557106 234178 557342 234414
rect 557426 234178 557662 234414
rect 557106 198498 557342 198734
rect 557426 198498 557662 198734
rect 557106 198178 557342 198414
rect 557426 198178 557662 198414
rect 557106 162498 557342 162734
rect 557426 162498 557662 162734
rect 557106 162178 557342 162414
rect 557426 162178 557662 162414
rect 557106 126498 557342 126734
rect 557426 126498 557662 126734
rect 557106 126178 557342 126414
rect 557426 126178 557662 126414
rect 557106 90498 557342 90734
rect 557426 90498 557662 90734
rect 557106 90178 557342 90414
rect 557426 90178 557662 90414
rect 557106 54498 557342 54734
rect 557426 54498 557662 54734
rect 557106 54178 557342 54414
rect 557426 54178 557662 54414
rect 557106 18498 557342 18734
rect 557426 18498 557662 18734
rect 557106 18178 557342 18414
rect 557426 18178 557662 18414
rect 557106 -4422 557342 -4186
rect 557426 -4422 557662 -4186
rect 557106 -4742 557342 -4506
rect 557426 -4742 557662 -4506
rect 560826 709402 561062 709638
rect 561146 709402 561382 709638
rect 560826 709082 561062 709318
rect 561146 709082 561382 709318
rect 560826 670218 561062 670454
rect 561146 670218 561382 670454
rect 560826 669898 561062 670134
rect 561146 669898 561382 670134
rect 560826 634218 561062 634454
rect 561146 634218 561382 634454
rect 560826 633898 561062 634134
rect 561146 633898 561382 634134
rect 560826 598218 561062 598454
rect 561146 598218 561382 598454
rect 560826 597898 561062 598134
rect 561146 597898 561382 598134
rect 560826 562218 561062 562454
rect 561146 562218 561382 562454
rect 560826 561898 561062 562134
rect 561146 561898 561382 562134
rect 560826 526218 561062 526454
rect 561146 526218 561382 526454
rect 560826 525898 561062 526134
rect 561146 525898 561382 526134
rect 560826 490218 561062 490454
rect 561146 490218 561382 490454
rect 560826 489898 561062 490134
rect 561146 489898 561382 490134
rect 560826 454218 561062 454454
rect 561146 454218 561382 454454
rect 560826 453898 561062 454134
rect 561146 453898 561382 454134
rect 560826 418218 561062 418454
rect 561146 418218 561382 418454
rect 560826 417898 561062 418134
rect 561146 417898 561382 418134
rect 560826 382218 561062 382454
rect 561146 382218 561382 382454
rect 560826 381898 561062 382134
rect 561146 381898 561382 382134
rect 560826 346218 561062 346454
rect 561146 346218 561382 346454
rect 560826 345898 561062 346134
rect 561146 345898 561382 346134
rect 560826 310218 561062 310454
rect 561146 310218 561382 310454
rect 560826 309898 561062 310134
rect 561146 309898 561382 310134
rect 560826 274218 561062 274454
rect 561146 274218 561382 274454
rect 560826 273898 561062 274134
rect 561146 273898 561382 274134
rect 560826 238218 561062 238454
rect 561146 238218 561382 238454
rect 560826 237898 561062 238134
rect 561146 237898 561382 238134
rect 560826 202218 561062 202454
rect 561146 202218 561382 202454
rect 560826 201898 561062 202134
rect 561146 201898 561382 202134
rect 560826 166218 561062 166454
rect 561146 166218 561382 166454
rect 560826 165898 561062 166134
rect 561146 165898 561382 166134
rect 560826 130218 561062 130454
rect 561146 130218 561382 130454
rect 560826 129898 561062 130134
rect 561146 129898 561382 130134
rect 560826 94218 561062 94454
rect 561146 94218 561382 94454
rect 560826 93898 561062 94134
rect 561146 93898 561382 94134
rect 560826 58218 561062 58454
rect 561146 58218 561382 58454
rect 560826 57898 561062 58134
rect 561146 57898 561382 58134
rect 560826 22218 561062 22454
rect 561146 22218 561382 22454
rect 560826 21898 561062 22134
rect 561146 21898 561382 22134
rect 560826 -5382 561062 -5146
rect 561146 -5382 561382 -5146
rect 560826 -5702 561062 -5466
rect 561146 -5702 561382 -5466
rect 564546 710362 564782 710598
rect 564866 710362 565102 710598
rect 564546 710042 564782 710278
rect 564866 710042 565102 710278
rect 564546 673938 564782 674174
rect 564866 673938 565102 674174
rect 564546 673618 564782 673854
rect 564866 673618 565102 673854
rect 564546 637938 564782 638174
rect 564866 637938 565102 638174
rect 564546 637618 564782 637854
rect 564866 637618 565102 637854
rect 564546 601938 564782 602174
rect 564866 601938 565102 602174
rect 564546 601618 564782 601854
rect 564866 601618 565102 601854
rect 564546 565938 564782 566174
rect 564866 565938 565102 566174
rect 564546 565618 564782 565854
rect 564866 565618 565102 565854
rect 564546 529938 564782 530174
rect 564866 529938 565102 530174
rect 564546 529618 564782 529854
rect 564866 529618 565102 529854
rect 564546 493938 564782 494174
rect 564866 493938 565102 494174
rect 564546 493618 564782 493854
rect 564866 493618 565102 493854
rect 564546 457938 564782 458174
rect 564866 457938 565102 458174
rect 564546 457618 564782 457854
rect 564866 457618 565102 457854
rect 564546 421938 564782 422174
rect 564866 421938 565102 422174
rect 564546 421618 564782 421854
rect 564866 421618 565102 421854
rect 564546 385938 564782 386174
rect 564866 385938 565102 386174
rect 564546 385618 564782 385854
rect 564866 385618 565102 385854
rect 564546 349938 564782 350174
rect 564866 349938 565102 350174
rect 564546 349618 564782 349854
rect 564866 349618 565102 349854
rect 564546 313938 564782 314174
rect 564866 313938 565102 314174
rect 564546 313618 564782 313854
rect 564866 313618 565102 313854
rect 564546 277938 564782 278174
rect 564866 277938 565102 278174
rect 564546 277618 564782 277854
rect 564866 277618 565102 277854
rect 564546 241938 564782 242174
rect 564866 241938 565102 242174
rect 564546 241618 564782 241854
rect 564866 241618 565102 241854
rect 564546 205938 564782 206174
rect 564866 205938 565102 206174
rect 564546 205618 564782 205854
rect 564866 205618 565102 205854
rect 564546 169938 564782 170174
rect 564866 169938 565102 170174
rect 564546 169618 564782 169854
rect 564866 169618 565102 169854
rect 564546 133938 564782 134174
rect 564866 133938 565102 134174
rect 564546 133618 564782 133854
rect 564866 133618 565102 133854
rect 564546 97938 564782 98174
rect 564866 97938 565102 98174
rect 564546 97618 564782 97854
rect 564866 97618 565102 97854
rect 564546 61938 564782 62174
rect 564866 61938 565102 62174
rect 564546 61618 564782 61854
rect 564866 61618 565102 61854
rect 564546 25938 564782 26174
rect 564866 25938 565102 26174
rect 564546 25618 564782 25854
rect 564866 25618 565102 25854
rect 564546 -6342 564782 -6106
rect 564866 -6342 565102 -6106
rect 564546 -6662 564782 -6426
rect 564866 -6662 565102 -6426
rect 568266 711322 568502 711558
rect 568586 711322 568822 711558
rect 568266 711002 568502 711238
rect 568586 711002 568822 711238
rect 568266 677658 568502 677894
rect 568586 677658 568822 677894
rect 568266 677338 568502 677574
rect 568586 677338 568822 677574
rect 568266 641658 568502 641894
rect 568586 641658 568822 641894
rect 568266 641338 568502 641574
rect 568586 641338 568822 641574
rect 568266 605658 568502 605894
rect 568586 605658 568822 605894
rect 568266 605338 568502 605574
rect 568586 605338 568822 605574
rect 568266 569658 568502 569894
rect 568586 569658 568822 569894
rect 568266 569338 568502 569574
rect 568586 569338 568822 569574
rect 568266 533658 568502 533894
rect 568586 533658 568822 533894
rect 568266 533338 568502 533574
rect 568586 533338 568822 533574
rect 568266 497658 568502 497894
rect 568586 497658 568822 497894
rect 568266 497338 568502 497574
rect 568586 497338 568822 497574
rect 568266 461658 568502 461894
rect 568586 461658 568822 461894
rect 568266 461338 568502 461574
rect 568586 461338 568822 461574
rect 568266 425658 568502 425894
rect 568586 425658 568822 425894
rect 568266 425338 568502 425574
rect 568586 425338 568822 425574
rect 568266 389658 568502 389894
rect 568586 389658 568822 389894
rect 568266 389338 568502 389574
rect 568586 389338 568822 389574
rect 568266 353658 568502 353894
rect 568586 353658 568822 353894
rect 568266 353338 568502 353574
rect 568586 353338 568822 353574
rect 568266 317658 568502 317894
rect 568586 317658 568822 317894
rect 568266 317338 568502 317574
rect 568586 317338 568822 317574
rect 568266 281658 568502 281894
rect 568586 281658 568822 281894
rect 568266 281338 568502 281574
rect 568586 281338 568822 281574
rect 568266 245658 568502 245894
rect 568586 245658 568822 245894
rect 568266 245338 568502 245574
rect 568586 245338 568822 245574
rect 568266 209658 568502 209894
rect 568586 209658 568822 209894
rect 568266 209338 568502 209574
rect 568586 209338 568822 209574
rect 568266 173658 568502 173894
rect 568586 173658 568822 173894
rect 568266 173338 568502 173574
rect 568586 173338 568822 173574
rect 568266 137658 568502 137894
rect 568586 137658 568822 137894
rect 568266 137338 568502 137574
rect 568586 137338 568822 137574
rect 568266 101658 568502 101894
rect 568586 101658 568822 101894
rect 568266 101338 568502 101574
rect 568586 101338 568822 101574
rect 568266 65658 568502 65894
rect 568586 65658 568822 65894
rect 568266 65338 568502 65574
rect 568586 65338 568822 65574
rect 568266 29658 568502 29894
rect 568586 29658 568822 29894
rect 568266 29338 568502 29574
rect 568586 29338 568822 29574
rect 568266 -7302 568502 -7066
rect 568586 -7302 568822 -7066
rect 568266 -7622 568502 -7386
rect 568586 -7622 568822 -7386
rect 578226 704602 578462 704838
rect 578546 704602 578782 704838
rect 578226 704282 578462 704518
rect 578546 704282 578782 704518
rect 578226 687618 578462 687854
rect 578546 687618 578782 687854
rect 578226 687298 578462 687534
rect 578546 687298 578782 687534
rect 578226 651618 578462 651854
rect 578546 651618 578782 651854
rect 578226 651298 578462 651534
rect 578546 651298 578782 651534
rect 578226 615618 578462 615854
rect 578546 615618 578782 615854
rect 578226 615298 578462 615534
rect 578546 615298 578782 615534
rect 578226 579618 578462 579854
rect 578546 579618 578782 579854
rect 578226 579298 578462 579534
rect 578546 579298 578782 579534
rect 578226 543618 578462 543854
rect 578546 543618 578782 543854
rect 578226 543298 578462 543534
rect 578546 543298 578782 543534
rect 578226 507618 578462 507854
rect 578546 507618 578782 507854
rect 578226 507298 578462 507534
rect 578546 507298 578782 507534
rect 578226 471618 578462 471854
rect 578546 471618 578782 471854
rect 578226 471298 578462 471534
rect 578546 471298 578782 471534
rect 578226 435618 578462 435854
rect 578546 435618 578782 435854
rect 578226 435298 578462 435534
rect 578546 435298 578782 435534
rect 578226 399618 578462 399854
rect 578546 399618 578782 399854
rect 578226 399298 578462 399534
rect 578546 399298 578782 399534
rect 578226 363618 578462 363854
rect 578546 363618 578782 363854
rect 578226 363298 578462 363534
rect 578546 363298 578782 363534
rect 578226 327618 578462 327854
rect 578546 327618 578782 327854
rect 578226 327298 578462 327534
rect 578546 327298 578782 327534
rect 578226 291618 578462 291854
rect 578546 291618 578782 291854
rect 578226 291298 578462 291534
rect 578546 291298 578782 291534
rect 578226 255618 578462 255854
rect 578546 255618 578782 255854
rect 578226 255298 578462 255534
rect 578546 255298 578782 255534
rect 578226 219618 578462 219854
rect 578546 219618 578782 219854
rect 578226 219298 578462 219534
rect 578546 219298 578782 219534
rect 578226 183618 578462 183854
rect 578546 183618 578782 183854
rect 578226 183298 578462 183534
rect 578546 183298 578782 183534
rect 578226 147618 578462 147854
rect 578546 147618 578782 147854
rect 578226 147298 578462 147534
rect 578546 147298 578782 147534
rect 578226 111618 578462 111854
rect 578546 111618 578782 111854
rect 578226 111298 578462 111534
rect 578546 111298 578782 111534
rect 578226 75618 578462 75854
rect 578546 75618 578782 75854
rect 578226 75298 578462 75534
rect 578546 75298 578782 75534
rect 578226 39618 578462 39854
rect 578546 39618 578782 39854
rect 578226 39298 578462 39534
rect 578546 39298 578782 39534
rect 578226 3618 578462 3854
rect 578546 3618 578782 3854
rect 578226 3298 578462 3534
rect 578546 3298 578782 3534
rect 578226 -582 578462 -346
rect 578546 -582 578782 -346
rect 578226 -902 578462 -666
rect 578546 -902 578782 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581946 705562 582182 705798
rect 582266 705562 582502 705798
rect 581946 705242 582182 705478
rect 582266 705242 582502 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581946 691338 582182 691574
rect 582266 691338 582502 691574
rect 581946 691018 582182 691254
rect 582266 691018 582502 691254
rect 581946 655338 582182 655574
rect 582266 655338 582502 655574
rect 581946 655018 582182 655254
rect 582266 655018 582502 655254
rect 581946 619338 582182 619574
rect 582266 619338 582502 619574
rect 581946 619018 582182 619254
rect 582266 619018 582502 619254
rect 581946 583338 582182 583574
rect 582266 583338 582502 583574
rect 581946 583018 582182 583254
rect 582266 583018 582502 583254
rect 581946 547338 582182 547574
rect 582266 547338 582502 547574
rect 581946 547018 582182 547254
rect 582266 547018 582502 547254
rect 581946 511338 582182 511574
rect 582266 511338 582502 511574
rect 581946 511018 582182 511254
rect 582266 511018 582502 511254
rect 581946 475338 582182 475574
rect 582266 475338 582502 475574
rect 581946 475018 582182 475254
rect 582266 475018 582502 475254
rect 581946 439338 582182 439574
rect 582266 439338 582502 439574
rect 581946 439018 582182 439254
rect 582266 439018 582502 439254
rect 581946 403338 582182 403574
rect 582266 403338 582502 403574
rect 581946 403018 582182 403254
rect 582266 403018 582502 403254
rect 581946 367338 582182 367574
rect 582266 367338 582502 367574
rect 581946 367018 582182 367254
rect 582266 367018 582502 367254
rect 581946 331338 582182 331574
rect 582266 331338 582502 331574
rect 581946 331018 582182 331254
rect 582266 331018 582502 331254
rect 581946 295338 582182 295574
rect 582266 295338 582502 295574
rect 581946 295018 582182 295254
rect 582266 295018 582502 295254
rect 581946 259338 582182 259574
rect 582266 259338 582502 259574
rect 581946 259018 582182 259254
rect 582266 259018 582502 259254
rect 581946 223338 582182 223574
rect 582266 223338 582502 223574
rect 581946 223018 582182 223254
rect 582266 223018 582502 223254
rect 581946 187338 582182 187574
rect 582266 187338 582502 187574
rect 581946 187018 582182 187254
rect 582266 187018 582502 187254
rect 581946 151338 582182 151574
rect 582266 151338 582502 151574
rect 581946 151018 582182 151254
rect 582266 151018 582502 151254
rect 581946 115338 582182 115574
rect 582266 115338 582502 115574
rect 581946 115018 582182 115254
rect 582266 115018 582502 115254
rect 581946 79338 582182 79574
rect 582266 79338 582502 79574
rect 581946 79018 582182 79254
rect 582266 79018 582502 79254
rect 581946 43338 582182 43574
rect 582266 43338 582502 43574
rect 581946 43018 582182 43254
rect 582266 43018 582502 43254
rect 581946 7338 582182 7574
rect 582266 7338 582502 7574
rect 581946 7018 582182 7254
rect 582266 7018 582502 7254
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687618 585578 687854
rect 585662 687618 585898 687854
rect 585342 687298 585578 687534
rect 585662 687298 585898 687534
rect 585342 651618 585578 651854
rect 585662 651618 585898 651854
rect 585342 651298 585578 651534
rect 585662 651298 585898 651534
rect 585342 615618 585578 615854
rect 585662 615618 585898 615854
rect 585342 615298 585578 615534
rect 585662 615298 585898 615534
rect 585342 579618 585578 579854
rect 585662 579618 585898 579854
rect 585342 579298 585578 579534
rect 585662 579298 585898 579534
rect 585342 543618 585578 543854
rect 585662 543618 585898 543854
rect 585342 543298 585578 543534
rect 585662 543298 585898 543534
rect 585342 507618 585578 507854
rect 585662 507618 585898 507854
rect 585342 507298 585578 507534
rect 585662 507298 585898 507534
rect 585342 471618 585578 471854
rect 585662 471618 585898 471854
rect 585342 471298 585578 471534
rect 585662 471298 585898 471534
rect 585342 435618 585578 435854
rect 585662 435618 585898 435854
rect 585342 435298 585578 435534
rect 585662 435298 585898 435534
rect 585342 399618 585578 399854
rect 585662 399618 585898 399854
rect 585342 399298 585578 399534
rect 585662 399298 585898 399534
rect 585342 363618 585578 363854
rect 585662 363618 585898 363854
rect 585342 363298 585578 363534
rect 585662 363298 585898 363534
rect 585342 327618 585578 327854
rect 585662 327618 585898 327854
rect 585342 327298 585578 327534
rect 585662 327298 585898 327534
rect 585342 291618 585578 291854
rect 585662 291618 585898 291854
rect 585342 291298 585578 291534
rect 585662 291298 585898 291534
rect 585342 255618 585578 255854
rect 585662 255618 585898 255854
rect 585342 255298 585578 255534
rect 585662 255298 585898 255534
rect 585342 219618 585578 219854
rect 585662 219618 585898 219854
rect 585342 219298 585578 219534
rect 585662 219298 585898 219534
rect 585342 183618 585578 183854
rect 585662 183618 585898 183854
rect 585342 183298 585578 183534
rect 585662 183298 585898 183534
rect 585342 147618 585578 147854
rect 585662 147618 585898 147854
rect 585342 147298 585578 147534
rect 585662 147298 585898 147534
rect 585342 111618 585578 111854
rect 585662 111618 585898 111854
rect 585342 111298 585578 111534
rect 585662 111298 585898 111534
rect 585342 75618 585578 75854
rect 585662 75618 585898 75854
rect 585342 75298 585578 75534
rect 585662 75298 585898 75534
rect 585342 39618 585578 39854
rect 585662 39618 585898 39854
rect 585342 39298 585578 39534
rect 585662 39298 585898 39534
rect 585342 3618 585578 3854
rect 585662 3618 585898 3854
rect 585342 3298 585578 3534
rect 585662 3298 585898 3534
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691338 586538 691574
rect 586622 691338 586858 691574
rect 586302 691018 586538 691254
rect 586622 691018 586858 691254
rect 586302 655338 586538 655574
rect 586622 655338 586858 655574
rect 586302 655018 586538 655254
rect 586622 655018 586858 655254
rect 586302 619338 586538 619574
rect 586622 619338 586858 619574
rect 586302 619018 586538 619254
rect 586622 619018 586858 619254
rect 586302 583338 586538 583574
rect 586622 583338 586858 583574
rect 586302 583018 586538 583254
rect 586622 583018 586858 583254
rect 586302 547338 586538 547574
rect 586622 547338 586858 547574
rect 586302 547018 586538 547254
rect 586622 547018 586858 547254
rect 586302 511338 586538 511574
rect 586622 511338 586858 511574
rect 586302 511018 586538 511254
rect 586622 511018 586858 511254
rect 586302 475338 586538 475574
rect 586622 475338 586858 475574
rect 586302 475018 586538 475254
rect 586622 475018 586858 475254
rect 586302 439338 586538 439574
rect 586622 439338 586858 439574
rect 586302 439018 586538 439254
rect 586622 439018 586858 439254
rect 586302 403338 586538 403574
rect 586622 403338 586858 403574
rect 586302 403018 586538 403254
rect 586622 403018 586858 403254
rect 586302 367338 586538 367574
rect 586622 367338 586858 367574
rect 586302 367018 586538 367254
rect 586622 367018 586858 367254
rect 586302 331338 586538 331574
rect 586622 331338 586858 331574
rect 586302 331018 586538 331254
rect 586622 331018 586858 331254
rect 586302 295338 586538 295574
rect 586622 295338 586858 295574
rect 586302 295018 586538 295254
rect 586622 295018 586858 295254
rect 586302 259338 586538 259574
rect 586622 259338 586858 259574
rect 586302 259018 586538 259254
rect 586622 259018 586858 259254
rect 586302 223338 586538 223574
rect 586622 223338 586858 223574
rect 586302 223018 586538 223254
rect 586622 223018 586858 223254
rect 586302 187338 586538 187574
rect 586622 187338 586858 187574
rect 586302 187018 586538 187254
rect 586622 187018 586858 187254
rect 586302 151338 586538 151574
rect 586622 151338 586858 151574
rect 586302 151018 586538 151254
rect 586622 151018 586858 151254
rect 586302 115338 586538 115574
rect 586622 115338 586858 115574
rect 586302 115018 586538 115254
rect 586622 115018 586858 115254
rect 586302 79338 586538 79574
rect 586622 79338 586858 79574
rect 586302 79018 586538 79254
rect 586622 79018 586858 79254
rect 586302 43338 586538 43574
rect 586622 43338 586858 43574
rect 586302 43018 586538 43254
rect 586622 43018 586858 43254
rect 586302 7338 586538 7574
rect 586622 7338 586858 7574
rect 586302 7018 586538 7254
rect 586622 7018 586858 7254
rect 581946 -1542 582182 -1306
rect 582266 -1542 582502 -1306
rect 581946 -1862 582182 -1626
rect 582266 -1862 582502 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 695058 587498 695294
rect 587582 695058 587818 695294
rect 587262 694738 587498 694974
rect 587582 694738 587818 694974
rect 587262 659058 587498 659294
rect 587582 659058 587818 659294
rect 587262 658738 587498 658974
rect 587582 658738 587818 658974
rect 587262 623058 587498 623294
rect 587582 623058 587818 623294
rect 587262 622738 587498 622974
rect 587582 622738 587818 622974
rect 587262 587058 587498 587294
rect 587582 587058 587818 587294
rect 587262 586738 587498 586974
rect 587582 586738 587818 586974
rect 587262 551058 587498 551294
rect 587582 551058 587818 551294
rect 587262 550738 587498 550974
rect 587582 550738 587818 550974
rect 587262 515058 587498 515294
rect 587582 515058 587818 515294
rect 587262 514738 587498 514974
rect 587582 514738 587818 514974
rect 587262 479058 587498 479294
rect 587582 479058 587818 479294
rect 587262 478738 587498 478974
rect 587582 478738 587818 478974
rect 587262 443058 587498 443294
rect 587582 443058 587818 443294
rect 587262 442738 587498 442974
rect 587582 442738 587818 442974
rect 587262 407058 587498 407294
rect 587582 407058 587818 407294
rect 587262 406738 587498 406974
rect 587582 406738 587818 406974
rect 587262 371058 587498 371294
rect 587582 371058 587818 371294
rect 587262 370738 587498 370974
rect 587582 370738 587818 370974
rect 587262 335058 587498 335294
rect 587582 335058 587818 335294
rect 587262 334738 587498 334974
rect 587582 334738 587818 334974
rect 587262 299058 587498 299294
rect 587582 299058 587818 299294
rect 587262 298738 587498 298974
rect 587582 298738 587818 298974
rect 587262 263058 587498 263294
rect 587582 263058 587818 263294
rect 587262 262738 587498 262974
rect 587582 262738 587818 262974
rect 587262 227058 587498 227294
rect 587582 227058 587818 227294
rect 587262 226738 587498 226974
rect 587582 226738 587818 226974
rect 587262 191058 587498 191294
rect 587582 191058 587818 191294
rect 587262 190738 587498 190974
rect 587582 190738 587818 190974
rect 587262 155058 587498 155294
rect 587582 155058 587818 155294
rect 587262 154738 587498 154974
rect 587582 154738 587818 154974
rect 587262 119058 587498 119294
rect 587582 119058 587818 119294
rect 587262 118738 587498 118974
rect 587582 118738 587818 118974
rect 587262 83058 587498 83294
rect 587582 83058 587818 83294
rect 587262 82738 587498 82974
rect 587582 82738 587818 82974
rect 587262 47058 587498 47294
rect 587582 47058 587818 47294
rect 587262 46738 587498 46974
rect 587582 46738 587818 46974
rect 587262 11058 587498 11294
rect 587582 11058 587818 11294
rect 587262 10738 587498 10974
rect 587582 10738 587818 10974
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698778 588458 699014
rect 588542 698778 588778 699014
rect 588222 698458 588458 698694
rect 588542 698458 588778 698694
rect 588222 662778 588458 663014
rect 588542 662778 588778 663014
rect 588222 662458 588458 662694
rect 588542 662458 588778 662694
rect 588222 626778 588458 627014
rect 588542 626778 588778 627014
rect 588222 626458 588458 626694
rect 588542 626458 588778 626694
rect 588222 590778 588458 591014
rect 588542 590778 588778 591014
rect 588222 590458 588458 590694
rect 588542 590458 588778 590694
rect 588222 554778 588458 555014
rect 588542 554778 588778 555014
rect 588222 554458 588458 554694
rect 588542 554458 588778 554694
rect 588222 518778 588458 519014
rect 588542 518778 588778 519014
rect 588222 518458 588458 518694
rect 588542 518458 588778 518694
rect 588222 482778 588458 483014
rect 588542 482778 588778 483014
rect 588222 482458 588458 482694
rect 588542 482458 588778 482694
rect 588222 446778 588458 447014
rect 588542 446778 588778 447014
rect 588222 446458 588458 446694
rect 588542 446458 588778 446694
rect 588222 410778 588458 411014
rect 588542 410778 588778 411014
rect 588222 410458 588458 410694
rect 588542 410458 588778 410694
rect 588222 374778 588458 375014
rect 588542 374778 588778 375014
rect 588222 374458 588458 374694
rect 588542 374458 588778 374694
rect 588222 338778 588458 339014
rect 588542 338778 588778 339014
rect 588222 338458 588458 338694
rect 588542 338458 588778 338694
rect 588222 302778 588458 303014
rect 588542 302778 588778 303014
rect 588222 302458 588458 302694
rect 588542 302458 588778 302694
rect 588222 266778 588458 267014
rect 588542 266778 588778 267014
rect 588222 266458 588458 266694
rect 588542 266458 588778 266694
rect 588222 230778 588458 231014
rect 588542 230778 588778 231014
rect 588222 230458 588458 230694
rect 588542 230458 588778 230694
rect 588222 194778 588458 195014
rect 588542 194778 588778 195014
rect 588222 194458 588458 194694
rect 588542 194458 588778 194694
rect 588222 158778 588458 159014
rect 588542 158778 588778 159014
rect 588222 158458 588458 158694
rect 588542 158458 588778 158694
rect 588222 122778 588458 123014
rect 588542 122778 588778 123014
rect 588222 122458 588458 122694
rect 588542 122458 588778 122694
rect 588222 86778 588458 87014
rect 588542 86778 588778 87014
rect 588222 86458 588458 86694
rect 588542 86458 588778 86694
rect 588222 50778 588458 51014
rect 588542 50778 588778 51014
rect 588222 50458 588458 50694
rect 588542 50458 588778 50694
rect 588222 14778 588458 15014
rect 588542 14778 588778 15014
rect 588222 14458 588458 14694
rect 588542 14458 588778 14694
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666498 589418 666734
rect 589502 666498 589738 666734
rect 589182 666178 589418 666414
rect 589502 666178 589738 666414
rect 589182 630498 589418 630734
rect 589502 630498 589738 630734
rect 589182 630178 589418 630414
rect 589502 630178 589738 630414
rect 589182 594498 589418 594734
rect 589502 594498 589738 594734
rect 589182 594178 589418 594414
rect 589502 594178 589738 594414
rect 589182 558498 589418 558734
rect 589502 558498 589738 558734
rect 589182 558178 589418 558414
rect 589502 558178 589738 558414
rect 589182 522498 589418 522734
rect 589502 522498 589738 522734
rect 589182 522178 589418 522414
rect 589502 522178 589738 522414
rect 589182 486498 589418 486734
rect 589502 486498 589738 486734
rect 589182 486178 589418 486414
rect 589502 486178 589738 486414
rect 589182 450498 589418 450734
rect 589502 450498 589738 450734
rect 589182 450178 589418 450414
rect 589502 450178 589738 450414
rect 589182 414498 589418 414734
rect 589502 414498 589738 414734
rect 589182 414178 589418 414414
rect 589502 414178 589738 414414
rect 589182 378498 589418 378734
rect 589502 378498 589738 378734
rect 589182 378178 589418 378414
rect 589502 378178 589738 378414
rect 589182 342498 589418 342734
rect 589502 342498 589738 342734
rect 589182 342178 589418 342414
rect 589502 342178 589738 342414
rect 589182 306498 589418 306734
rect 589502 306498 589738 306734
rect 589182 306178 589418 306414
rect 589502 306178 589738 306414
rect 589182 270498 589418 270734
rect 589502 270498 589738 270734
rect 589182 270178 589418 270414
rect 589502 270178 589738 270414
rect 589182 234498 589418 234734
rect 589502 234498 589738 234734
rect 589182 234178 589418 234414
rect 589502 234178 589738 234414
rect 589182 198498 589418 198734
rect 589502 198498 589738 198734
rect 589182 198178 589418 198414
rect 589502 198178 589738 198414
rect 589182 162498 589418 162734
rect 589502 162498 589738 162734
rect 589182 162178 589418 162414
rect 589502 162178 589738 162414
rect 589182 126498 589418 126734
rect 589502 126498 589738 126734
rect 589182 126178 589418 126414
rect 589502 126178 589738 126414
rect 589182 90498 589418 90734
rect 589502 90498 589738 90734
rect 589182 90178 589418 90414
rect 589502 90178 589738 90414
rect 589182 54498 589418 54734
rect 589502 54498 589738 54734
rect 589182 54178 589418 54414
rect 589502 54178 589738 54414
rect 589182 18498 589418 18734
rect 589502 18498 589738 18734
rect 589182 18178 589418 18414
rect 589502 18178 589738 18414
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 670218 590378 670454
rect 590462 670218 590698 670454
rect 590142 669898 590378 670134
rect 590462 669898 590698 670134
rect 590142 634218 590378 634454
rect 590462 634218 590698 634454
rect 590142 633898 590378 634134
rect 590462 633898 590698 634134
rect 590142 598218 590378 598454
rect 590462 598218 590698 598454
rect 590142 597898 590378 598134
rect 590462 597898 590698 598134
rect 590142 562218 590378 562454
rect 590462 562218 590698 562454
rect 590142 561898 590378 562134
rect 590462 561898 590698 562134
rect 590142 526218 590378 526454
rect 590462 526218 590698 526454
rect 590142 525898 590378 526134
rect 590462 525898 590698 526134
rect 590142 490218 590378 490454
rect 590462 490218 590698 490454
rect 590142 489898 590378 490134
rect 590462 489898 590698 490134
rect 590142 454218 590378 454454
rect 590462 454218 590698 454454
rect 590142 453898 590378 454134
rect 590462 453898 590698 454134
rect 590142 418218 590378 418454
rect 590462 418218 590698 418454
rect 590142 417898 590378 418134
rect 590462 417898 590698 418134
rect 590142 382218 590378 382454
rect 590462 382218 590698 382454
rect 590142 381898 590378 382134
rect 590462 381898 590698 382134
rect 590142 346218 590378 346454
rect 590462 346218 590698 346454
rect 590142 345898 590378 346134
rect 590462 345898 590698 346134
rect 590142 310218 590378 310454
rect 590462 310218 590698 310454
rect 590142 309898 590378 310134
rect 590462 309898 590698 310134
rect 590142 274218 590378 274454
rect 590462 274218 590698 274454
rect 590142 273898 590378 274134
rect 590462 273898 590698 274134
rect 590142 238218 590378 238454
rect 590462 238218 590698 238454
rect 590142 237898 590378 238134
rect 590462 237898 590698 238134
rect 590142 202218 590378 202454
rect 590462 202218 590698 202454
rect 590142 201898 590378 202134
rect 590462 201898 590698 202134
rect 590142 166218 590378 166454
rect 590462 166218 590698 166454
rect 590142 165898 590378 166134
rect 590462 165898 590698 166134
rect 590142 130218 590378 130454
rect 590462 130218 590698 130454
rect 590142 129898 590378 130134
rect 590462 129898 590698 130134
rect 590142 94218 590378 94454
rect 590462 94218 590698 94454
rect 590142 93898 590378 94134
rect 590462 93898 590698 94134
rect 590142 58218 590378 58454
rect 590462 58218 590698 58454
rect 590142 57898 590378 58134
rect 590462 57898 590698 58134
rect 590142 22218 590378 22454
rect 590462 22218 590698 22454
rect 590142 21898 590378 22134
rect 590462 21898 590698 22134
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673938 591338 674174
rect 591422 673938 591658 674174
rect 591102 673618 591338 673854
rect 591422 673618 591658 673854
rect 591102 637938 591338 638174
rect 591422 637938 591658 638174
rect 591102 637618 591338 637854
rect 591422 637618 591658 637854
rect 591102 601938 591338 602174
rect 591422 601938 591658 602174
rect 591102 601618 591338 601854
rect 591422 601618 591658 601854
rect 591102 565938 591338 566174
rect 591422 565938 591658 566174
rect 591102 565618 591338 565854
rect 591422 565618 591658 565854
rect 591102 529938 591338 530174
rect 591422 529938 591658 530174
rect 591102 529618 591338 529854
rect 591422 529618 591658 529854
rect 591102 493938 591338 494174
rect 591422 493938 591658 494174
rect 591102 493618 591338 493854
rect 591422 493618 591658 493854
rect 591102 457938 591338 458174
rect 591422 457938 591658 458174
rect 591102 457618 591338 457854
rect 591422 457618 591658 457854
rect 591102 421938 591338 422174
rect 591422 421938 591658 422174
rect 591102 421618 591338 421854
rect 591422 421618 591658 421854
rect 591102 385938 591338 386174
rect 591422 385938 591658 386174
rect 591102 385618 591338 385854
rect 591422 385618 591658 385854
rect 591102 349938 591338 350174
rect 591422 349938 591658 350174
rect 591102 349618 591338 349854
rect 591422 349618 591658 349854
rect 591102 313938 591338 314174
rect 591422 313938 591658 314174
rect 591102 313618 591338 313854
rect 591422 313618 591658 313854
rect 591102 277938 591338 278174
rect 591422 277938 591658 278174
rect 591102 277618 591338 277854
rect 591422 277618 591658 277854
rect 591102 241938 591338 242174
rect 591422 241938 591658 242174
rect 591102 241618 591338 241854
rect 591422 241618 591658 241854
rect 591102 205938 591338 206174
rect 591422 205938 591658 206174
rect 591102 205618 591338 205854
rect 591422 205618 591658 205854
rect 591102 169938 591338 170174
rect 591422 169938 591658 170174
rect 591102 169618 591338 169854
rect 591422 169618 591658 169854
rect 591102 133938 591338 134174
rect 591422 133938 591658 134174
rect 591102 133618 591338 133854
rect 591422 133618 591658 133854
rect 591102 97938 591338 98174
rect 591422 97938 591658 98174
rect 591102 97618 591338 97854
rect 591422 97618 591658 97854
rect 591102 61938 591338 62174
rect 591422 61938 591658 62174
rect 591102 61618 591338 61854
rect 591422 61618 591658 61854
rect 591102 25938 591338 26174
rect 591422 25938 591658 26174
rect 591102 25618 591338 25854
rect 591422 25618 591658 25854
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677658 592298 677894
rect 592382 677658 592618 677894
rect 592062 677338 592298 677574
rect 592382 677338 592618 677574
rect 592062 641658 592298 641894
rect 592382 641658 592618 641894
rect 592062 641338 592298 641574
rect 592382 641338 592618 641574
rect 592062 605658 592298 605894
rect 592382 605658 592618 605894
rect 592062 605338 592298 605574
rect 592382 605338 592618 605574
rect 592062 569658 592298 569894
rect 592382 569658 592618 569894
rect 592062 569338 592298 569574
rect 592382 569338 592618 569574
rect 592062 533658 592298 533894
rect 592382 533658 592618 533894
rect 592062 533338 592298 533574
rect 592382 533338 592618 533574
rect 592062 497658 592298 497894
rect 592382 497658 592618 497894
rect 592062 497338 592298 497574
rect 592382 497338 592618 497574
rect 592062 461658 592298 461894
rect 592382 461658 592618 461894
rect 592062 461338 592298 461574
rect 592382 461338 592618 461574
rect 592062 425658 592298 425894
rect 592382 425658 592618 425894
rect 592062 425338 592298 425574
rect 592382 425338 592618 425574
rect 592062 389658 592298 389894
rect 592382 389658 592618 389894
rect 592062 389338 592298 389574
rect 592382 389338 592618 389574
rect 592062 353658 592298 353894
rect 592382 353658 592618 353894
rect 592062 353338 592298 353574
rect 592382 353338 592618 353574
rect 592062 317658 592298 317894
rect 592382 317658 592618 317894
rect 592062 317338 592298 317574
rect 592382 317338 592618 317574
rect 592062 281658 592298 281894
rect 592382 281658 592618 281894
rect 592062 281338 592298 281574
rect 592382 281338 592618 281574
rect 592062 245658 592298 245894
rect 592382 245658 592618 245894
rect 592062 245338 592298 245574
rect 592382 245338 592618 245574
rect 592062 209658 592298 209894
rect 592382 209658 592618 209894
rect 592062 209338 592298 209574
rect 592382 209338 592618 209574
rect 592062 173658 592298 173894
rect 592382 173658 592618 173894
rect 592062 173338 592298 173574
rect 592382 173338 592618 173574
rect 592062 137658 592298 137894
rect 592382 137658 592618 137894
rect 592062 137338 592298 137574
rect 592382 137338 592618 137574
rect 592062 101658 592298 101894
rect 592382 101658 592618 101894
rect 592062 101338 592298 101574
rect 592382 101338 592618 101574
rect 592062 65658 592298 65894
rect 592382 65658 592618 65894
rect 592062 65338 592298 65574
rect 592382 65338 592618 65574
rect 592062 29658 592298 29894
rect 592382 29658 592618 29894
rect 592062 29338 592298 29574
rect 592382 29338 592618 29574
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 28266 711558
rect 28502 711322 28586 711558
rect 28822 711322 64266 711558
rect 64502 711322 64586 711558
rect 64822 711322 100266 711558
rect 100502 711322 100586 711558
rect 100822 711322 136266 711558
rect 136502 711322 136586 711558
rect 136822 711322 172266 711558
rect 172502 711322 172586 711558
rect 172822 711322 208266 711558
rect 208502 711322 208586 711558
rect 208822 711322 244266 711558
rect 244502 711322 244586 711558
rect 244822 711322 280266 711558
rect 280502 711322 280586 711558
rect 280822 711322 316266 711558
rect 316502 711322 316586 711558
rect 316822 711322 352266 711558
rect 352502 711322 352586 711558
rect 352822 711322 388266 711558
rect 388502 711322 388586 711558
rect 388822 711322 424266 711558
rect 424502 711322 424586 711558
rect 424822 711322 460266 711558
rect 460502 711322 460586 711558
rect 460822 711322 496266 711558
rect 496502 711322 496586 711558
rect 496822 711322 532266 711558
rect 532502 711322 532586 711558
rect 532822 711322 568266 711558
rect 568502 711322 568586 711558
rect 568822 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 28266 711238
rect 28502 711002 28586 711238
rect 28822 711002 64266 711238
rect 64502 711002 64586 711238
rect 64822 711002 100266 711238
rect 100502 711002 100586 711238
rect 100822 711002 136266 711238
rect 136502 711002 136586 711238
rect 136822 711002 172266 711238
rect 172502 711002 172586 711238
rect 172822 711002 208266 711238
rect 208502 711002 208586 711238
rect 208822 711002 244266 711238
rect 244502 711002 244586 711238
rect 244822 711002 280266 711238
rect 280502 711002 280586 711238
rect 280822 711002 316266 711238
rect 316502 711002 316586 711238
rect 316822 711002 352266 711238
rect 352502 711002 352586 711238
rect 352822 711002 388266 711238
rect 388502 711002 388586 711238
rect 388822 711002 424266 711238
rect 424502 711002 424586 711238
rect 424822 711002 460266 711238
rect 460502 711002 460586 711238
rect 460822 711002 496266 711238
rect 496502 711002 496586 711238
rect 496822 711002 532266 711238
rect 532502 711002 532586 711238
rect 532822 711002 568266 711238
rect 568502 711002 568586 711238
rect 568822 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24546 710598
rect 24782 710362 24866 710598
rect 25102 710362 60546 710598
rect 60782 710362 60866 710598
rect 61102 710362 96546 710598
rect 96782 710362 96866 710598
rect 97102 710362 132546 710598
rect 132782 710362 132866 710598
rect 133102 710362 168546 710598
rect 168782 710362 168866 710598
rect 169102 710362 204546 710598
rect 204782 710362 204866 710598
rect 205102 710362 240546 710598
rect 240782 710362 240866 710598
rect 241102 710362 276546 710598
rect 276782 710362 276866 710598
rect 277102 710362 312546 710598
rect 312782 710362 312866 710598
rect 313102 710362 348546 710598
rect 348782 710362 348866 710598
rect 349102 710362 384546 710598
rect 384782 710362 384866 710598
rect 385102 710362 420546 710598
rect 420782 710362 420866 710598
rect 421102 710362 456546 710598
rect 456782 710362 456866 710598
rect 457102 710362 492546 710598
rect 492782 710362 492866 710598
rect 493102 710362 528546 710598
rect 528782 710362 528866 710598
rect 529102 710362 564546 710598
rect 564782 710362 564866 710598
rect 565102 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24546 710278
rect 24782 710042 24866 710278
rect 25102 710042 60546 710278
rect 60782 710042 60866 710278
rect 61102 710042 96546 710278
rect 96782 710042 96866 710278
rect 97102 710042 132546 710278
rect 132782 710042 132866 710278
rect 133102 710042 168546 710278
rect 168782 710042 168866 710278
rect 169102 710042 204546 710278
rect 204782 710042 204866 710278
rect 205102 710042 240546 710278
rect 240782 710042 240866 710278
rect 241102 710042 276546 710278
rect 276782 710042 276866 710278
rect 277102 710042 312546 710278
rect 312782 710042 312866 710278
rect 313102 710042 348546 710278
rect 348782 710042 348866 710278
rect 349102 710042 384546 710278
rect 384782 710042 384866 710278
rect 385102 710042 420546 710278
rect 420782 710042 420866 710278
rect 421102 710042 456546 710278
rect 456782 710042 456866 710278
rect 457102 710042 492546 710278
rect 492782 710042 492866 710278
rect 493102 710042 528546 710278
rect 528782 710042 528866 710278
rect 529102 710042 564546 710278
rect 564782 710042 564866 710278
rect 565102 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20826 709638
rect 21062 709402 21146 709638
rect 21382 709402 56826 709638
rect 57062 709402 57146 709638
rect 57382 709402 92826 709638
rect 93062 709402 93146 709638
rect 93382 709402 128826 709638
rect 129062 709402 129146 709638
rect 129382 709402 164826 709638
rect 165062 709402 165146 709638
rect 165382 709402 200826 709638
rect 201062 709402 201146 709638
rect 201382 709402 236826 709638
rect 237062 709402 237146 709638
rect 237382 709402 272826 709638
rect 273062 709402 273146 709638
rect 273382 709402 308826 709638
rect 309062 709402 309146 709638
rect 309382 709402 344826 709638
rect 345062 709402 345146 709638
rect 345382 709402 380826 709638
rect 381062 709402 381146 709638
rect 381382 709402 416826 709638
rect 417062 709402 417146 709638
rect 417382 709402 452826 709638
rect 453062 709402 453146 709638
rect 453382 709402 488826 709638
rect 489062 709402 489146 709638
rect 489382 709402 524826 709638
rect 525062 709402 525146 709638
rect 525382 709402 560826 709638
rect 561062 709402 561146 709638
rect 561382 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20826 709318
rect 21062 709082 21146 709318
rect 21382 709082 56826 709318
rect 57062 709082 57146 709318
rect 57382 709082 92826 709318
rect 93062 709082 93146 709318
rect 93382 709082 128826 709318
rect 129062 709082 129146 709318
rect 129382 709082 164826 709318
rect 165062 709082 165146 709318
rect 165382 709082 200826 709318
rect 201062 709082 201146 709318
rect 201382 709082 236826 709318
rect 237062 709082 237146 709318
rect 237382 709082 272826 709318
rect 273062 709082 273146 709318
rect 273382 709082 308826 709318
rect 309062 709082 309146 709318
rect 309382 709082 344826 709318
rect 345062 709082 345146 709318
rect 345382 709082 380826 709318
rect 381062 709082 381146 709318
rect 381382 709082 416826 709318
rect 417062 709082 417146 709318
rect 417382 709082 452826 709318
rect 453062 709082 453146 709318
rect 453382 709082 488826 709318
rect 489062 709082 489146 709318
rect 489382 709082 524826 709318
rect 525062 709082 525146 709318
rect 525382 709082 560826 709318
rect 561062 709082 561146 709318
rect 561382 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 17106 708678
rect 17342 708442 17426 708678
rect 17662 708442 53106 708678
rect 53342 708442 53426 708678
rect 53662 708442 89106 708678
rect 89342 708442 89426 708678
rect 89662 708442 125106 708678
rect 125342 708442 125426 708678
rect 125662 708442 161106 708678
rect 161342 708442 161426 708678
rect 161662 708442 197106 708678
rect 197342 708442 197426 708678
rect 197662 708442 233106 708678
rect 233342 708442 233426 708678
rect 233662 708442 269106 708678
rect 269342 708442 269426 708678
rect 269662 708442 305106 708678
rect 305342 708442 305426 708678
rect 305662 708442 341106 708678
rect 341342 708442 341426 708678
rect 341662 708442 377106 708678
rect 377342 708442 377426 708678
rect 377662 708442 413106 708678
rect 413342 708442 413426 708678
rect 413662 708442 449106 708678
rect 449342 708442 449426 708678
rect 449662 708442 485106 708678
rect 485342 708442 485426 708678
rect 485662 708442 521106 708678
rect 521342 708442 521426 708678
rect 521662 708442 557106 708678
rect 557342 708442 557426 708678
rect 557662 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 17106 708358
rect 17342 708122 17426 708358
rect 17662 708122 53106 708358
rect 53342 708122 53426 708358
rect 53662 708122 89106 708358
rect 89342 708122 89426 708358
rect 89662 708122 125106 708358
rect 125342 708122 125426 708358
rect 125662 708122 161106 708358
rect 161342 708122 161426 708358
rect 161662 708122 197106 708358
rect 197342 708122 197426 708358
rect 197662 708122 233106 708358
rect 233342 708122 233426 708358
rect 233662 708122 269106 708358
rect 269342 708122 269426 708358
rect 269662 708122 305106 708358
rect 305342 708122 305426 708358
rect 305662 708122 341106 708358
rect 341342 708122 341426 708358
rect 341662 708122 377106 708358
rect 377342 708122 377426 708358
rect 377662 708122 413106 708358
rect 413342 708122 413426 708358
rect 413662 708122 449106 708358
rect 449342 708122 449426 708358
rect 449662 708122 485106 708358
rect 485342 708122 485426 708358
rect 485662 708122 521106 708358
rect 521342 708122 521426 708358
rect 521662 708122 557106 708358
rect 557342 708122 557426 708358
rect 557662 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 13386 707718
rect 13622 707482 13706 707718
rect 13942 707482 49386 707718
rect 49622 707482 49706 707718
rect 49942 707482 85386 707718
rect 85622 707482 85706 707718
rect 85942 707482 121386 707718
rect 121622 707482 121706 707718
rect 121942 707482 157386 707718
rect 157622 707482 157706 707718
rect 157942 707482 193386 707718
rect 193622 707482 193706 707718
rect 193942 707482 229386 707718
rect 229622 707482 229706 707718
rect 229942 707482 265386 707718
rect 265622 707482 265706 707718
rect 265942 707482 301386 707718
rect 301622 707482 301706 707718
rect 301942 707482 337386 707718
rect 337622 707482 337706 707718
rect 337942 707482 373386 707718
rect 373622 707482 373706 707718
rect 373942 707482 409386 707718
rect 409622 707482 409706 707718
rect 409942 707482 445386 707718
rect 445622 707482 445706 707718
rect 445942 707482 481386 707718
rect 481622 707482 481706 707718
rect 481942 707482 517386 707718
rect 517622 707482 517706 707718
rect 517942 707482 553386 707718
rect 553622 707482 553706 707718
rect 553942 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 13386 707398
rect 13622 707162 13706 707398
rect 13942 707162 49386 707398
rect 49622 707162 49706 707398
rect 49942 707162 85386 707398
rect 85622 707162 85706 707398
rect 85942 707162 121386 707398
rect 121622 707162 121706 707398
rect 121942 707162 157386 707398
rect 157622 707162 157706 707398
rect 157942 707162 193386 707398
rect 193622 707162 193706 707398
rect 193942 707162 229386 707398
rect 229622 707162 229706 707398
rect 229942 707162 265386 707398
rect 265622 707162 265706 707398
rect 265942 707162 301386 707398
rect 301622 707162 301706 707398
rect 301942 707162 337386 707398
rect 337622 707162 337706 707398
rect 337942 707162 373386 707398
rect 373622 707162 373706 707398
rect 373942 707162 409386 707398
rect 409622 707162 409706 707398
rect 409942 707162 445386 707398
rect 445622 707162 445706 707398
rect 445942 707162 481386 707398
rect 481622 707162 481706 707398
rect 481942 707162 517386 707398
rect 517622 707162 517706 707398
rect 517942 707162 553386 707398
rect 553622 707162 553706 707398
rect 553942 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9666 706758
rect 9902 706522 9986 706758
rect 10222 706522 45666 706758
rect 45902 706522 45986 706758
rect 46222 706522 81666 706758
rect 81902 706522 81986 706758
rect 82222 706522 117666 706758
rect 117902 706522 117986 706758
rect 118222 706522 153666 706758
rect 153902 706522 153986 706758
rect 154222 706522 189666 706758
rect 189902 706522 189986 706758
rect 190222 706522 225666 706758
rect 225902 706522 225986 706758
rect 226222 706522 261666 706758
rect 261902 706522 261986 706758
rect 262222 706522 297666 706758
rect 297902 706522 297986 706758
rect 298222 706522 333666 706758
rect 333902 706522 333986 706758
rect 334222 706522 369666 706758
rect 369902 706522 369986 706758
rect 370222 706522 405666 706758
rect 405902 706522 405986 706758
rect 406222 706522 441666 706758
rect 441902 706522 441986 706758
rect 442222 706522 477666 706758
rect 477902 706522 477986 706758
rect 478222 706522 513666 706758
rect 513902 706522 513986 706758
rect 514222 706522 549666 706758
rect 549902 706522 549986 706758
rect 550222 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9666 706438
rect 9902 706202 9986 706438
rect 10222 706202 45666 706438
rect 45902 706202 45986 706438
rect 46222 706202 81666 706438
rect 81902 706202 81986 706438
rect 82222 706202 117666 706438
rect 117902 706202 117986 706438
rect 118222 706202 153666 706438
rect 153902 706202 153986 706438
rect 154222 706202 189666 706438
rect 189902 706202 189986 706438
rect 190222 706202 225666 706438
rect 225902 706202 225986 706438
rect 226222 706202 261666 706438
rect 261902 706202 261986 706438
rect 262222 706202 297666 706438
rect 297902 706202 297986 706438
rect 298222 706202 333666 706438
rect 333902 706202 333986 706438
rect 334222 706202 369666 706438
rect 369902 706202 369986 706438
rect 370222 706202 405666 706438
rect 405902 706202 405986 706438
rect 406222 706202 441666 706438
rect 441902 706202 441986 706438
rect 442222 706202 477666 706438
rect 477902 706202 477986 706438
rect 478222 706202 513666 706438
rect 513902 706202 513986 706438
rect 514222 706202 549666 706438
rect 549902 706202 549986 706438
rect 550222 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5946 705798
rect 6182 705562 6266 705798
rect 6502 705562 41946 705798
rect 42182 705562 42266 705798
rect 42502 705562 77946 705798
rect 78182 705562 78266 705798
rect 78502 705562 113946 705798
rect 114182 705562 114266 705798
rect 114502 705562 149946 705798
rect 150182 705562 150266 705798
rect 150502 705562 185946 705798
rect 186182 705562 186266 705798
rect 186502 705562 221946 705798
rect 222182 705562 222266 705798
rect 222502 705562 257946 705798
rect 258182 705562 258266 705798
rect 258502 705562 293946 705798
rect 294182 705562 294266 705798
rect 294502 705562 329946 705798
rect 330182 705562 330266 705798
rect 330502 705562 365946 705798
rect 366182 705562 366266 705798
rect 366502 705562 401946 705798
rect 402182 705562 402266 705798
rect 402502 705562 437946 705798
rect 438182 705562 438266 705798
rect 438502 705562 473946 705798
rect 474182 705562 474266 705798
rect 474502 705562 509946 705798
rect 510182 705562 510266 705798
rect 510502 705562 545946 705798
rect 546182 705562 546266 705798
rect 546502 705562 581946 705798
rect 582182 705562 582266 705798
rect 582502 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5946 705478
rect 6182 705242 6266 705478
rect 6502 705242 41946 705478
rect 42182 705242 42266 705478
rect 42502 705242 77946 705478
rect 78182 705242 78266 705478
rect 78502 705242 113946 705478
rect 114182 705242 114266 705478
rect 114502 705242 149946 705478
rect 150182 705242 150266 705478
rect 150502 705242 185946 705478
rect 186182 705242 186266 705478
rect 186502 705242 221946 705478
rect 222182 705242 222266 705478
rect 222502 705242 257946 705478
rect 258182 705242 258266 705478
rect 258502 705242 293946 705478
rect 294182 705242 294266 705478
rect 294502 705242 329946 705478
rect 330182 705242 330266 705478
rect 330502 705242 365946 705478
rect 366182 705242 366266 705478
rect 366502 705242 401946 705478
rect 402182 705242 402266 705478
rect 402502 705242 437946 705478
rect 438182 705242 438266 705478
rect 438502 705242 473946 705478
rect 474182 705242 474266 705478
rect 474502 705242 509946 705478
rect 510182 705242 510266 705478
rect 510502 705242 545946 705478
rect 546182 705242 546266 705478
rect 546502 705242 581946 705478
rect 582182 705242 582266 705478
rect 582502 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 2226 704838
rect 2462 704602 2546 704838
rect 2782 704602 38226 704838
rect 38462 704602 38546 704838
rect 38782 704602 74226 704838
rect 74462 704602 74546 704838
rect 74782 704602 110226 704838
rect 110462 704602 110546 704838
rect 110782 704602 146226 704838
rect 146462 704602 146546 704838
rect 146782 704602 182226 704838
rect 182462 704602 182546 704838
rect 182782 704602 218226 704838
rect 218462 704602 218546 704838
rect 218782 704602 254226 704838
rect 254462 704602 254546 704838
rect 254782 704602 290226 704838
rect 290462 704602 290546 704838
rect 290782 704602 326226 704838
rect 326462 704602 326546 704838
rect 326782 704602 362226 704838
rect 362462 704602 362546 704838
rect 362782 704602 398226 704838
rect 398462 704602 398546 704838
rect 398782 704602 434226 704838
rect 434462 704602 434546 704838
rect 434782 704602 470226 704838
rect 470462 704602 470546 704838
rect 470782 704602 506226 704838
rect 506462 704602 506546 704838
rect 506782 704602 542226 704838
rect 542462 704602 542546 704838
rect 542782 704602 578226 704838
rect 578462 704602 578546 704838
rect 578782 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 2226 704518
rect 2462 704282 2546 704518
rect 2782 704282 38226 704518
rect 38462 704282 38546 704518
rect 38782 704282 74226 704518
rect 74462 704282 74546 704518
rect 74782 704282 110226 704518
rect 110462 704282 110546 704518
rect 110782 704282 146226 704518
rect 146462 704282 146546 704518
rect 146782 704282 182226 704518
rect 182462 704282 182546 704518
rect 182782 704282 218226 704518
rect 218462 704282 218546 704518
rect 218782 704282 254226 704518
rect 254462 704282 254546 704518
rect 254782 704282 290226 704518
rect 290462 704282 290546 704518
rect 290782 704282 326226 704518
rect 326462 704282 326546 704518
rect 326782 704282 362226 704518
rect 362462 704282 362546 704518
rect 362782 704282 398226 704518
rect 398462 704282 398546 704518
rect 398782 704282 434226 704518
rect 434462 704282 434546 704518
rect 434782 704282 470226 704518
rect 470462 704282 470546 704518
rect 470782 704282 506226 704518
rect 506462 704282 506546 704518
rect 506782 704282 542226 704518
rect 542462 704282 542546 704518
rect 542782 704282 578226 704518
rect 578462 704282 578546 704518
rect 578782 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 699014 592650 699046
rect -8726 698778 -4854 699014
rect -4618 698778 -4534 699014
rect -4298 698778 13386 699014
rect 13622 698778 13706 699014
rect 13942 698778 49386 699014
rect 49622 698778 49706 699014
rect 49942 698778 85386 699014
rect 85622 698778 85706 699014
rect 85942 698778 121386 699014
rect 121622 698778 121706 699014
rect 121942 698778 157386 699014
rect 157622 698778 157706 699014
rect 157942 698778 193386 699014
rect 193622 698778 193706 699014
rect 193942 698778 229386 699014
rect 229622 698778 229706 699014
rect 229942 698778 265386 699014
rect 265622 698778 265706 699014
rect 265942 698778 301386 699014
rect 301622 698778 301706 699014
rect 301942 698778 337386 699014
rect 337622 698778 337706 699014
rect 337942 698778 373386 699014
rect 373622 698778 373706 699014
rect 373942 698778 409386 699014
rect 409622 698778 409706 699014
rect 409942 698778 445386 699014
rect 445622 698778 445706 699014
rect 445942 698778 481386 699014
rect 481622 698778 481706 699014
rect 481942 698778 517386 699014
rect 517622 698778 517706 699014
rect 517942 698778 553386 699014
rect 553622 698778 553706 699014
rect 553942 698778 588222 699014
rect 588458 698778 588542 699014
rect 588778 698778 592650 699014
rect -8726 698694 592650 698778
rect -8726 698458 -4854 698694
rect -4618 698458 -4534 698694
rect -4298 698458 13386 698694
rect 13622 698458 13706 698694
rect 13942 698458 49386 698694
rect 49622 698458 49706 698694
rect 49942 698458 85386 698694
rect 85622 698458 85706 698694
rect 85942 698458 121386 698694
rect 121622 698458 121706 698694
rect 121942 698458 157386 698694
rect 157622 698458 157706 698694
rect 157942 698458 193386 698694
rect 193622 698458 193706 698694
rect 193942 698458 229386 698694
rect 229622 698458 229706 698694
rect 229942 698458 265386 698694
rect 265622 698458 265706 698694
rect 265942 698458 301386 698694
rect 301622 698458 301706 698694
rect 301942 698458 337386 698694
rect 337622 698458 337706 698694
rect 337942 698458 373386 698694
rect 373622 698458 373706 698694
rect 373942 698458 409386 698694
rect 409622 698458 409706 698694
rect 409942 698458 445386 698694
rect 445622 698458 445706 698694
rect 445942 698458 481386 698694
rect 481622 698458 481706 698694
rect 481942 698458 517386 698694
rect 517622 698458 517706 698694
rect 517942 698458 553386 698694
rect 553622 698458 553706 698694
rect 553942 698458 588222 698694
rect 588458 698458 588542 698694
rect 588778 698458 592650 698694
rect -8726 698426 592650 698458
rect -8726 695294 592650 695326
rect -8726 695058 -3894 695294
rect -3658 695058 -3574 695294
rect -3338 695058 9666 695294
rect 9902 695058 9986 695294
rect 10222 695058 45666 695294
rect 45902 695058 45986 695294
rect 46222 695058 81666 695294
rect 81902 695058 81986 695294
rect 82222 695058 117666 695294
rect 117902 695058 117986 695294
rect 118222 695058 153666 695294
rect 153902 695058 153986 695294
rect 154222 695058 189666 695294
rect 189902 695058 189986 695294
rect 190222 695058 225666 695294
rect 225902 695058 225986 695294
rect 226222 695058 261666 695294
rect 261902 695058 261986 695294
rect 262222 695058 297666 695294
rect 297902 695058 297986 695294
rect 298222 695058 333666 695294
rect 333902 695058 333986 695294
rect 334222 695058 369666 695294
rect 369902 695058 369986 695294
rect 370222 695058 405666 695294
rect 405902 695058 405986 695294
rect 406222 695058 441666 695294
rect 441902 695058 441986 695294
rect 442222 695058 477666 695294
rect 477902 695058 477986 695294
rect 478222 695058 513666 695294
rect 513902 695058 513986 695294
rect 514222 695058 549666 695294
rect 549902 695058 549986 695294
rect 550222 695058 587262 695294
rect 587498 695058 587582 695294
rect 587818 695058 592650 695294
rect -8726 694974 592650 695058
rect -8726 694738 -3894 694974
rect -3658 694738 -3574 694974
rect -3338 694738 9666 694974
rect 9902 694738 9986 694974
rect 10222 694738 45666 694974
rect 45902 694738 45986 694974
rect 46222 694738 81666 694974
rect 81902 694738 81986 694974
rect 82222 694738 117666 694974
rect 117902 694738 117986 694974
rect 118222 694738 153666 694974
rect 153902 694738 153986 694974
rect 154222 694738 189666 694974
rect 189902 694738 189986 694974
rect 190222 694738 225666 694974
rect 225902 694738 225986 694974
rect 226222 694738 261666 694974
rect 261902 694738 261986 694974
rect 262222 694738 297666 694974
rect 297902 694738 297986 694974
rect 298222 694738 333666 694974
rect 333902 694738 333986 694974
rect 334222 694738 369666 694974
rect 369902 694738 369986 694974
rect 370222 694738 405666 694974
rect 405902 694738 405986 694974
rect 406222 694738 441666 694974
rect 441902 694738 441986 694974
rect 442222 694738 477666 694974
rect 477902 694738 477986 694974
rect 478222 694738 513666 694974
rect 513902 694738 513986 694974
rect 514222 694738 549666 694974
rect 549902 694738 549986 694974
rect 550222 694738 587262 694974
rect 587498 694738 587582 694974
rect 587818 694738 592650 694974
rect -8726 694706 592650 694738
rect -8726 691574 592650 691606
rect -8726 691338 -2934 691574
rect -2698 691338 -2614 691574
rect -2378 691338 5946 691574
rect 6182 691338 6266 691574
rect 6502 691338 41946 691574
rect 42182 691338 42266 691574
rect 42502 691338 77946 691574
rect 78182 691338 78266 691574
rect 78502 691338 113946 691574
rect 114182 691338 114266 691574
rect 114502 691338 149946 691574
rect 150182 691338 150266 691574
rect 150502 691338 185946 691574
rect 186182 691338 186266 691574
rect 186502 691338 221946 691574
rect 222182 691338 222266 691574
rect 222502 691338 257946 691574
rect 258182 691338 258266 691574
rect 258502 691338 293946 691574
rect 294182 691338 294266 691574
rect 294502 691338 329946 691574
rect 330182 691338 330266 691574
rect 330502 691338 365946 691574
rect 366182 691338 366266 691574
rect 366502 691338 401946 691574
rect 402182 691338 402266 691574
rect 402502 691338 437946 691574
rect 438182 691338 438266 691574
rect 438502 691338 473946 691574
rect 474182 691338 474266 691574
rect 474502 691338 509946 691574
rect 510182 691338 510266 691574
rect 510502 691338 545946 691574
rect 546182 691338 546266 691574
rect 546502 691338 581946 691574
rect 582182 691338 582266 691574
rect 582502 691338 586302 691574
rect 586538 691338 586622 691574
rect 586858 691338 592650 691574
rect -8726 691254 592650 691338
rect -8726 691018 -2934 691254
rect -2698 691018 -2614 691254
rect -2378 691018 5946 691254
rect 6182 691018 6266 691254
rect 6502 691018 41946 691254
rect 42182 691018 42266 691254
rect 42502 691018 77946 691254
rect 78182 691018 78266 691254
rect 78502 691018 113946 691254
rect 114182 691018 114266 691254
rect 114502 691018 149946 691254
rect 150182 691018 150266 691254
rect 150502 691018 185946 691254
rect 186182 691018 186266 691254
rect 186502 691018 221946 691254
rect 222182 691018 222266 691254
rect 222502 691018 257946 691254
rect 258182 691018 258266 691254
rect 258502 691018 293946 691254
rect 294182 691018 294266 691254
rect 294502 691018 329946 691254
rect 330182 691018 330266 691254
rect 330502 691018 365946 691254
rect 366182 691018 366266 691254
rect 366502 691018 401946 691254
rect 402182 691018 402266 691254
rect 402502 691018 437946 691254
rect 438182 691018 438266 691254
rect 438502 691018 473946 691254
rect 474182 691018 474266 691254
rect 474502 691018 509946 691254
rect 510182 691018 510266 691254
rect 510502 691018 545946 691254
rect 546182 691018 546266 691254
rect 546502 691018 581946 691254
rect 582182 691018 582266 691254
rect 582502 691018 586302 691254
rect 586538 691018 586622 691254
rect 586858 691018 592650 691254
rect -8726 690986 592650 691018
rect -8726 687854 592650 687886
rect -8726 687618 -1974 687854
rect -1738 687618 -1654 687854
rect -1418 687618 2226 687854
rect 2462 687618 2546 687854
rect 2782 687618 38226 687854
rect 38462 687618 38546 687854
rect 38782 687618 74226 687854
rect 74462 687618 74546 687854
rect 74782 687618 110226 687854
rect 110462 687618 110546 687854
rect 110782 687618 146226 687854
rect 146462 687618 146546 687854
rect 146782 687618 182226 687854
rect 182462 687618 182546 687854
rect 182782 687618 218226 687854
rect 218462 687618 218546 687854
rect 218782 687618 254226 687854
rect 254462 687618 254546 687854
rect 254782 687618 290226 687854
rect 290462 687618 290546 687854
rect 290782 687618 326226 687854
rect 326462 687618 326546 687854
rect 326782 687618 362226 687854
rect 362462 687618 362546 687854
rect 362782 687618 398226 687854
rect 398462 687618 398546 687854
rect 398782 687618 434226 687854
rect 434462 687618 434546 687854
rect 434782 687618 470226 687854
rect 470462 687618 470546 687854
rect 470782 687618 506226 687854
rect 506462 687618 506546 687854
rect 506782 687618 542226 687854
rect 542462 687618 542546 687854
rect 542782 687618 578226 687854
rect 578462 687618 578546 687854
rect 578782 687618 585342 687854
rect 585578 687618 585662 687854
rect 585898 687618 592650 687854
rect -8726 687534 592650 687618
rect -8726 687298 -1974 687534
rect -1738 687298 -1654 687534
rect -1418 687298 2226 687534
rect 2462 687298 2546 687534
rect 2782 687298 38226 687534
rect 38462 687298 38546 687534
rect 38782 687298 74226 687534
rect 74462 687298 74546 687534
rect 74782 687298 110226 687534
rect 110462 687298 110546 687534
rect 110782 687298 146226 687534
rect 146462 687298 146546 687534
rect 146782 687298 182226 687534
rect 182462 687298 182546 687534
rect 182782 687298 218226 687534
rect 218462 687298 218546 687534
rect 218782 687298 254226 687534
rect 254462 687298 254546 687534
rect 254782 687298 290226 687534
rect 290462 687298 290546 687534
rect 290782 687298 326226 687534
rect 326462 687298 326546 687534
rect 326782 687298 362226 687534
rect 362462 687298 362546 687534
rect 362782 687298 398226 687534
rect 398462 687298 398546 687534
rect 398782 687298 434226 687534
rect 434462 687298 434546 687534
rect 434782 687298 470226 687534
rect 470462 687298 470546 687534
rect 470782 687298 506226 687534
rect 506462 687298 506546 687534
rect 506782 687298 542226 687534
rect 542462 687298 542546 687534
rect 542782 687298 578226 687534
rect 578462 687298 578546 687534
rect 578782 687298 585342 687534
rect 585578 687298 585662 687534
rect 585898 687298 592650 687534
rect -8726 687266 592650 687298
rect -8726 677894 592650 677926
rect -8726 677658 -8694 677894
rect -8458 677658 -8374 677894
rect -8138 677658 28266 677894
rect 28502 677658 28586 677894
rect 28822 677658 64266 677894
rect 64502 677658 64586 677894
rect 64822 677658 100266 677894
rect 100502 677658 100586 677894
rect 100822 677658 136266 677894
rect 136502 677658 136586 677894
rect 136822 677658 172266 677894
rect 172502 677658 172586 677894
rect 172822 677658 208266 677894
rect 208502 677658 208586 677894
rect 208822 677658 244266 677894
rect 244502 677658 244586 677894
rect 244822 677658 280266 677894
rect 280502 677658 280586 677894
rect 280822 677658 316266 677894
rect 316502 677658 316586 677894
rect 316822 677658 352266 677894
rect 352502 677658 352586 677894
rect 352822 677658 388266 677894
rect 388502 677658 388586 677894
rect 388822 677658 424266 677894
rect 424502 677658 424586 677894
rect 424822 677658 460266 677894
rect 460502 677658 460586 677894
rect 460822 677658 496266 677894
rect 496502 677658 496586 677894
rect 496822 677658 532266 677894
rect 532502 677658 532586 677894
rect 532822 677658 568266 677894
rect 568502 677658 568586 677894
rect 568822 677658 592062 677894
rect 592298 677658 592382 677894
rect 592618 677658 592650 677894
rect -8726 677574 592650 677658
rect -8726 677338 -8694 677574
rect -8458 677338 -8374 677574
rect -8138 677338 28266 677574
rect 28502 677338 28586 677574
rect 28822 677338 64266 677574
rect 64502 677338 64586 677574
rect 64822 677338 100266 677574
rect 100502 677338 100586 677574
rect 100822 677338 136266 677574
rect 136502 677338 136586 677574
rect 136822 677338 172266 677574
rect 172502 677338 172586 677574
rect 172822 677338 208266 677574
rect 208502 677338 208586 677574
rect 208822 677338 244266 677574
rect 244502 677338 244586 677574
rect 244822 677338 280266 677574
rect 280502 677338 280586 677574
rect 280822 677338 316266 677574
rect 316502 677338 316586 677574
rect 316822 677338 352266 677574
rect 352502 677338 352586 677574
rect 352822 677338 388266 677574
rect 388502 677338 388586 677574
rect 388822 677338 424266 677574
rect 424502 677338 424586 677574
rect 424822 677338 460266 677574
rect 460502 677338 460586 677574
rect 460822 677338 496266 677574
rect 496502 677338 496586 677574
rect 496822 677338 532266 677574
rect 532502 677338 532586 677574
rect 532822 677338 568266 677574
rect 568502 677338 568586 677574
rect 568822 677338 592062 677574
rect 592298 677338 592382 677574
rect 592618 677338 592650 677574
rect -8726 677306 592650 677338
rect -8726 674174 592650 674206
rect -8726 673938 -7734 674174
rect -7498 673938 -7414 674174
rect -7178 673938 24546 674174
rect 24782 673938 24866 674174
rect 25102 673938 60546 674174
rect 60782 673938 60866 674174
rect 61102 673938 96546 674174
rect 96782 673938 96866 674174
rect 97102 673938 132546 674174
rect 132782 673938 132866 674174
rect 133102 673938 168546 674174
rect 168782 673938 168866 674174
rect 169102 673938 204546 674174
rect 204782 673938 204866 674174
rect 205102 673938 240546 674174
rect 240782 673938 240866 674174
rect 241102 673938 276546 674174
rect 276782 673938 276866 674174
rect 277102 673938 312546 674174
rect 312782 673938 312866 674174
rect 313102 673938 348546 674174
rect 348782 673938 348866 674174
rect 349102 673938 384546 674174
rect 384782 673938 384866 674174
rect 385102 673938 420546 674174
rect 420782 673938 420866 674174
rect 421102 673938 456546 674174
rect 456782 673938 456866 674174
rect 457102 673938 492546 674174
rect 492782 673938 492866 674174
rect 493102 673938 528546 674174
rect 528782 673938 528866 674174
rect 529102 673938 564546 674174
rect 564782 673938 564866 674174
rect 565102 673938 591102 674174
rect 591338 673938 591422 674174
rect 591658 673938 592650 674174
rect -8726 673854 592650 673938
rect -8726 673618 -7734 673854
rect -7498 673618 -7414 673854
rect -7178 673618 24546 673854
rect 24782 673618 24866 673854
rect 25102 673618 60546 673854
rect 60782 673618 60866 673854
rect 61102 673618 96546 673854
rect 96782 673618 96866 673854
rect 97102 673618 132546 673854
rect 132782 673618 132866 673854
rect 133102 673618 168546 673854
rect 168782 673618 168866 673854
rect 169102 673618 204546 673854
rect 204782 673618 204866 673854
rect 205102 673618 240546 673854
rect 240782 673618 240866 673854
rect 241102 673618 276546 673854
rect 276782 673618 276866 673854
rect 277102 673618 312546 673854
rect 312782 673618 312866 673854
rect 313102 673618 348546 673854
rect 348782 673618 348866 673854
rect 349102 673618 384546 673854
rect 384782 673618 384866 673854
rect 385102 673618 420546 673854
rect 420782 673618 420866 673854
rect 421102 673618 456546 673854
rect 456782 673618 456866 673854
rect 457102 673618 492546 673854
rect 492782 673618 492866 673854
rect 493102 673618 528546 673854
rect 528782 673618 528866 673854
rect 529102 673618 564546 673854
rect 564782 673618 564866 673854
rect 565102 673618 591102 673854
rect 591338 673618 591422 673854
rect 591658 673618 592650 673854
rect -8726 673586 592650 673618
rect -8726 670454 592650 670486
rect -8726 670218 -6774 670454
rect -6538 670218 -6454 670454
rect -6218 670218 20826 670454
rect 21062 670218 21146 670454
rect 21382 670218 56826 670454
rect 57062 670218 57146 670454
rect 57382 670218 92826 670454
rect 93062 670218 93146 670454
rect 93382 670218 128826 670454
rect 129062 670218 129146 670454
rect 129382 670218 164826 670454
rect 165062 670218 165146 670454
rect 165382 670218 200826 670454
rect 201062 670218 201146 670454
rect 201382 670218 236826 670454
rect 237062 670218 237146 670454
rect 237382 670218 272826 670454
rect 273062 670218 273146 670454
rect 273382 670218 308826 670454
rect 309062 670218 309146 670454
rect 309382 670218 344826 670454
rect 345062 670218 345146 670454
rect 345382 670218 380826 670454
rect 381062 670218 381146 670454
rect 381382 670218 416826 670454
rect 417062 670218 417146 670454
rect 417382 670218 452826 670454
rect 453062 670218 453146 670454
rect 453382 670218 488826 670454
rect 489062 670218 489146 670454
rect 489382 670218 524826 670454
rect 525062 670218 525146 670454
rect 525382 670218 560826 670454
rect 561062 670218 561146 670454
rect 561382 670218 590142 670454
rect 590378 670218 590462 670454
rect 590698 670218 592650 670454
rect -8726 670134 592650 670218
rect -8726 669898 -6774 670134
rect -6538 669898 -6454 670134
rect -6218 669898 20826 670134
rect 21062 669898 21146 670134
rect 21382 669898 56826 670134
rect 57062 669898 57146 670134
rect 57382 669898 92826 670134
rect 93062 669898 93146 670134
rect 93382 669898 128826 670134
rect 129062 669898 129146 670134
rect 129382 669898 164826 670134
rect 165062 669898 165146 670134
rect 165382 669898 200826 670134
rect 201062 669898 201146 670134
rect 201382 669898 236826 670134
rect 237062 669898 237146 670134
rect 237382 669898 272826 670134
rect 273062 669898 273146 670134
rect 273382 669898 308826 670134
rect 309062 669898 309146 670134
rect 309382 669898 344826 670134
rect 345062 669898 345146 670134
rect 345382 669898 380826 670134
rect 381062 669898 381146 670134
rect 381382 669898 416826 670134
rect 417062 669898 417146 670134
rect 417382 669898 452826 670134
rect 453062 669898 453146 670134
rect 453382 669898 488826 670134
rect 489062 669898 489146 670134
rect 489382 669898 524826 670134
rect 525062 669898 525146 670134
rect 525382 669898 560826 670134
rect 561062 669898 561146 670134
rect 561382 669898 590142 670134
rect 590378 669898 590462 670134
rect 590698 669898 592650 670134
rect -8726 669866 592650 669898
rect -8726 666734 592650 666766
rect -8726 666498 -5814 666734
rect -5578 666498 -5494 666734
rect -5258 666498 17106 666734
rect 17342 666498 17426 666734
rect 17662 666498 53106 666734
rect 53342 666498 53426 666734
rect 53662 666498 89106 666734
rect 89342 666498 89426 666734
rect 89662 666498 125106 666734
rect 125342 666498 125426 666734
rect 125662 666498 161106 666734
rect 161342 666498 161426 666734
rect 161662 666498 197106 666734
rect 197342 666498 197426 666734
rect 197662 666498 233106 666734
rect 233342 666498 233426 666734
rect 233662 666498 269106 666734
rect 269342 666498 269426 666734
rect 269662 666498 305106 666734
rect 305342 666498 305426 666734
rect 305662 666498 341106 666734
rect 341342 666498 341426 666734
rect 341662 666498 377106 666734
rect 377342 666498 377426 666734
rect 377662 666498 413106 666734
rect 413342 666498 413426 666734
rect 413662 666498 449106 666734
rect 449342 666498 449426 666734
rect 449662 666498 485106 666734
rect 485342 666498 485426 666734
rect 485662 666498 521106 666734
rect 521342 666498 521426 666734
rect 521662 666498 557106 666734
rect 557342 666498 557426 666734
rect 557662 666498 589182 666734
rect 589418 666498 589502 666734
rect 589738 666498 592650 666734
rect -8726 666414 592650 666498
rect -8726 666178 -5814 666414
rect -5578 666178 -5494 666414
rect -5258 666178 17106 666414
rect 17342 666178 17426 666414
rect 17662 666178 53106 666414
rect 53342 666178 53426 666414
rect 53662 666178 89106 666414
rect 89342 666178 89426 666414
rect 89662 666178 125106 666414
rect 125342 666178 125426 666414
rect 125662 666178 161106 666414
rect 161342 666178 161426 666414
rect 161662 666178 197106 666414
rect 197342 666178 197426 666414
rect 197662 666178 233106 666414
rect 233342 666178 233426 666414
rect 233662 666178 269106 666414
rect 269342 666178 269426 666414
rect 269662 666178 305106 666414
rect 305342 666178 305426 666414
rect 305662 666178 341106 666414
rect 341342 666178 341426 666414
rect 341662 666178 377106 666414
rect 377342 666178 377426 666414
rect 377662 666178 413106 666414
rect 413342 666178 413426 666414
rect 413662 666178 449106 666414
rect 449342 666178 449426 666414
rect 449662 666178 485106 666414
rect 485342 666178 485426 666414
rect 485662 666178 521106 666414
rect 521342 666178 521426 666414
rect 521662 666178 557106 666414
rect 557342 666178 557426 666414
rect 557662 666178 589182 666414
rect 589418 666178 589502 666414
rect 589738 666178 592650 666414
rect -8726 666146 592650 666178
rect -8726 663014 592650 663046
rect -8726 662778 -4854 663014
rect -4618 662778 -4534 663014
rect -4298 662778 13386 663014
rect 13622 662778 13706 663014
rect 13942 662778 49386 663014
rect 49622 662778 49706 663014
rect 49942 662778 85386 663014
rect 85622 662778 85706 663014
rect 85942 662778 121386 663014
rect 121622 662778 121706 663014
rect 121942 662778 157386 663014
rect 157622 662778 157706 663014
rect 157942 662778 193386 663014
rect 193622 662778 193706 663014
rect 193942 662778 229386 663014
rect 229622 662778 229706 663014
rect 229942 662778 265386 663014
rect 265622 662778 265706 663014
rect 265942 662778 301386 663014
rect 301622 662778 301706 663014
rect 301942 662778 337386 663014
rect 337622 662778 337706 663014
rect 337942 662778 373386 663014
rect 373622 662778 373706 663014
rect 373942 662778 409386 663014
rect 409622 662778 409706 663014
rect 409942 662778 445386 663014
rect 445622 662778 445706 663014
rect 445942 662778 481386 663014
rect 481622 662778 481706 663014
rect 481942 662778 517386 663014
rect 517622 662778 517706 663014
rect 517942 662778 553386 663014
rect 553622 662778 553706 663014
rect 553942 662778 588222 663014
rect 588458 662778 588542 663014
rect 588778 662778 592650 663014
rect -8726 662694 592650 662778
rect -8726 662458 -4854 662694
rect -4618 662458 -4534 662694
rect -4298 662458 13386 662694
rect 13622 662458 13706 662694
rect 13942 662458 49386 662694
rect 49622 662458 49706 662694
rect 49942 662458 85386 662694
rect 85622 662458 85706 662694
rect 85942 662458 121386 662694
rect 121622 662458 121706 662694
rect 121942 662458 157386 662694
rect 157622 662458 157706 662694
rect 157942 662458 193386 662694
rect 193622 662458 193706 662694
rect 193942 662458 229386 662694
rect 229622 662458 229706 662694
rect 229942 662458 265386 662694
rect 265622 662458 265706 662694
rect 265942 662458 301386 662694
rect 301622 662458 301706 662694
rect 301942 662458 337386 662694
rect 337622 662458 337706 662694
rect 337942 662458 373386 662694
rect 373622 662458 373706 662694
rect 373942 662458 409386 662694
rect 409622 662458 409706 662694
rect 409942 662458 445386 662694
rect 445622 662458 445706 662694
rect 445942 662458 481386 662694
rect 481622 662458 481706 662694
rect 481942 662458 517386 662694
rect 517622 662458 517706 662694
rect 517942 662458 553386 662694
rect 553622 662458 553706 662694
rect 553942 662458 588222 662694
rect 588458 662458 588542 662694
rect 588778 662458 592650 662694
rect -8726 662426 592650 662458
rect -8726 659294 592650 659326
rect -8726 659058 -3894 659294
rect -3658 659058 -3574 659294
rect -3338 659058 9666 659294
rect 9902 659058 9986 659294
rect 10222 659058 45666 659294
rect 45902 659058 45986 659294
rect 46222 659058 81666 659294
rect 81902 659058 81986 659294
rect 82222 659058 117666 659294
rect 117902 659058 117986 659294
rect 118222 659058 153666 659294
rect 153902 659058 153986 659294
rect 154222 659058 189666 659294
rect 189902 659058 189986 659294
rect 190222 659058 225666 659294
rect 225902 659058 225986 659294
rect 226222 659058 261666 659294
rect 261902 659058 261986 659294
rect 262222 659058 297666 659294
rect 297902 659058 297986 659294
rect 298222 659058 333666 659294
rect 333902 659058 333986 659294
rect 334222 659058 369666 659294
rect 369902 659058 369986 659294
rect 370222 659058 405666 659294
rect 405902 659058 405986 659294
rect 406222 659058 441666 659294
rect 441902 659058 441986 659294
rect 442222 659058 477666 659294
rect 477902 659058 477986 659294
rect 478222 659058 513666 659294
rect 513902 659058 513986 659294
rect 514222 659058 549666 659294
rect 549902 659058 549986 659294
rect 550222 659058 587262 659294
rect 587498 659058 587582 659294
rect 587818 659058 592650 659294
rect -8726 658974 592650 659058
rect -8726 658738 -3894 658974
rect -3658 658738 -3574 658974
rect -3338 658738 9666 658974
rect 9902 658738 9986 658974
rect 10222 658738 45666 658974
rect 45902 658738 45986 658974
rect 46222 658738 81666 658974
rect 81902 658738 81986 658974
rect 82222 658738 117666 658974
rect 117902 658738 117986 658974
rect 118222 658738 153666 658974
rect 153902 658738 153986 658974
rect 154222 658738 189666 658974
rect 189902 658738 189986 658974
rect 190222 658738 225666 658974
rect 225902 658738 225986 658974
rect 226222 658738 261666 658974
rect 261902 658738 261986 658974
rect 262222 658738 297666 658974
rect 297902 658738 297986 658974
rect 298222 658738 333666 658974
rect 333902 658738 333986 658974
rect 334222 658738 369666 658974
rect 369902 658738 369986 658974
rect 370222 658738 405666 658974
rect 405902 658738 405986 658974
rect 406222 658738 441666 658974
rect 441902 658738 441986 658974
rect 442222 658738 477666 658974
rect 477902 658738 477986 658974
rect 478222 658738 513666 658974
rect 513902 658738 513986 658974
rect 514222 658738 549666 658974
rect 549902 658738 549986 658974
rect 550222 658738 587262 658974
rect 587498 658738 587582 658974
rect 587818 658738 592650 658974
rect -8726 658706 592650 658738
rect -8726 655574 592650 655606
rect -8726 655338 -2934 655574
rect -2698 655338 -2614 655574
rect -2378 655338 5946 655574
rect 6182 655338 6266 655574
rect 6502 655338 41946 655574
rect 42182 655338 42266 655574
rect 42502 655338 77946 655574
rect 78182 655338 78266 655574
rect 78502 655338 113946 655574
rect 114182 655338 114266 655574
rect 114502 655338 149946 655574
rect 150182 655338 150266 655574
rect 150502 655338 185946 655574
rect 186182 655338 186266 655574
rect 186502 655338 221946 655574
rect 222182 655338 222266 655574
rect 222502 655338 257946 655574
rect 258182 655338 258266 655574
rect 258502 655338 293946 655574
rect 294182 655338 294266 655574
rect 294502 655338 329946 655574
rect 330182 655338 330266 655574
rect 330502 655338 365946 655574
rect 366182 655338 366266 655574
rect 366502 655338 401946 655574
rect 402182 655338 402266 655574
rect 402502 655338 437946 655574
rect 438182 655338 438266 655574
rect 438502 655338 473946 655574
rect 474182 655338 474266 655574
rect 474502 655338 509946 655574
rect 510182 655338 510266 655574
rect 510502 655338 545946 655574
rect 546182 655338 546266 655574
rect 546502 655338 581946 655574
rect 582182 655338 582266 655574
rect 582502 655338 586302 655574
rect 586538 655338 586622 655574
rect 586858 655338 592650 655574
rect -8726 655254 592650 655338
rect -8726 655018 -2934 655254
rect -2698 655018 -2614 655254
rect -2378 655018 5946 655254
rect 6182 655018 6266 655254
rect 6502 655018 41946 655254
rect 42182 655018 42266 655254
rect 42502 655018 77946 655254
rect 78182 655018 78266 655254
rect 78502 655018 113946 655254
rect 114182 655018 114266 655254
rect 114502 655018 149946 655254
rect 150182 655018 150266 655254
rect 150502 655018 185946 655254
rect 186182 655018 186266 655254
rect 186502 655018 221946 655254
rect 222182 655018 222266 655254
rect 222502 655018 257946 655254
rect 258182 655018 258266 655254
rect 258502 655018 293946 655254
rect 294182 655018 294266 655254
rect 294502 655018 329946 655254
rect 330182 655018 330266 655254
rect 330502 655018 365946 655254
rect 366182 655018 366266 655254
rect 366502 655018 401946 655254
rect 402182 655018 402266 655254
rect 402502 655018 437946 655254
rect 438182 655018 438266 655254
rect 438502 655018 473946 655254
rect 474182 655018 474266 655254
rect 474502 655018 509946 655254
rect 510182 655018 510266 655254
rect 510502 655018 545946 655254
rect 546182 655018 546266 655254
rect 546502 655018 581946 655254
rect 582182 655018 582266 655254
rect 582502 655018 586302 655254
rect 586538 655018 586622 655254
rect 586858 655018 592650 655254
rect -8726 654986 592650 655018
rect -8726 651854 592650 651886
rect -8726 651618 -1974 651854
rect -1738 651618 -1654 651854
rect -1418 651618 2226 651854
rect 2462 651618 2546 651854
rect 2782 651618 38226 651854
rect 38462 651618 38546 651854
rect 38782 651618 74226 651854
rect 74462 651618 74546 651854
rect 74782 651618 110226 651854
rect 110462 651618 110546 651854
rect 110782 651618 146226 651854
rect 146462 651618 146546 651854
rect 146782 651618 182226 651854
rect 182462 651618 182546 651854
rect 182782 651618 218226 651854
rect 218462 651618 218546 651854
rect 218782 651618 254226 651854
rect 254462 651618 254546 651854
rect 254782 651618 290226 651854
rect 290462 651618 290546 651854
rect 290782 651618 326226 651854
rect 326462 651618 326546 651854
rect 326782 651618 362226 651854
rect 362462 651618 362546 651854
rect 362782 651618 398226 651854
rect 398462 651618 398546 651854
rect 398782 651618 434226 651854
rect 434462 651618 434546 651854
rect 434782 651618 470226 651854
rect 470462 651618 470546 651854
rect 470782 651618 506226 651854
rect 506462 651618 506546 651854
rect 506782 651618 542226 651854
rect 542462 651618 542546 651854
rect 542782 651618 578226 651854
rect 578462 651618 578546 651854
rect 578782 651618 585342 651854
rect 585578 651618 585662 651854
rect 585898 651618 592650 651854
rect -8726 651534 592650 651618
rect -8726 651298 -1974 651534
rect -1738 651298 -1654 651534
rect -1418 651298 2226 651534
rect 2462 651298 2546 651534
rect 2782 651298 38226 651534
rect 38462 651298 38546 651534
rect 38782 651298 74226 651534
rect 74462 651298 74546 651534
rect 74782 651298 110226 651534
rect 110462 651298 110546 651534
rect 110782 651298 146226 651534
rect 146462 651298 146546 651534
rect 146782 651298 182226 651534
rect 182462 651298 182546 651534
rect 182782 651298 218226 651534
rect 218462 651298 218546 651534
rect 218782 651298 254226 651534
rect 254462 651298 254546 651534
rect 254782 651298 290226 651534
rect 290462 651298 290546 651534
rect 290782 651298 326226 651534
rect 326462 651298 326546 651534
rect 326782 651298 362226 651534
rect 362462 651298 362546 651534
rect 362782 651298 398226 651534
rect 398462 651298 398546 651534
rect 398782 651298 434226 651534
rect 434462 651298 434546 651534
rect 434782 651298 470226 651534
rect 470462 651298 470546 651534
rect 470782 651298 506226 651534
rect 506462 651298 506546 651534
rect 506782 651298 542226 651534
rect 542462 651298 542546 651534
rect 542782 651298 578226 651534
rect 578462 651298 578546 651534
rect 578782 651298 585342 651534
rect 585578 651298 585662 651534
rect 585898 651298 592650 651534
rect -8726 651266 592650 651298
rect -8726 641894 592650 641926
rect -8726 641658 -8694 641894
rect -8458 641658 -8374 641894
rect -8138 641658 28266 641894
rect 28502 641658 28586 641894
rect 28822 641658 64266 641894
rect 64502 641658 64586 641894
rect 64822 641658 100266 641894
rect 100502 641658 100586 641894
rect 100822 641658 136266 641894
rect 136502 641658 136586 641894
rect 136822 641658 172266 641894
rect 172502 641658 172586 641894
rect 172822 641658 208266 641894
rect 208502 641658 208586 641894
rect 208822 641658 244266 641894
rect 244502 641658 244586 641894
rect 244822 641658 280266 641894
rect 280502 641658 280586 641894
rect 280822 641658 316266 641894
rect 316502 641658 316586 641894
rect 316822 641658 352266 641894
rect 352502 641658 352586 641894
rect 352822 641658 388266 641894
rect 388502 641658 388586 641894
rect 388822 641658 424266 641894
rect 424502 641658 424586 641894
rect 424822 641658 460266 641894
rect 460502 641658 460586 641894
rect 460822 641658 496266 641894
rect 496502 641658 496586 641894
rect 496822 641658 532266 641894
rect 532502 641658 532586 641894
rect 532822 641658 568266 641894
rect 568502 641658 568586 641894
rect 568822 641658 592062 641894
rect 592298 641658 592382 641894
rect 592618 641658 592650 641894
rect -8726 641574 592650 641658
rect -8726 641338 -8694 641574
rect -8458 641338 -8374 641574
rect -8138 641338 28266 641574
rect 28502 641338 28586 641574
rect 28822 641338 64266 641574
rect 64502 641338 64586 641574
rect 64822 641338 100266 641574
rect 100502 641338 100586 641574
rect 100822 641338 136266 641574
rect 136502 641338 136586 641574
rect 136822 641338 172266 641574
rect 172502 641338 172586 641574
rect 172822 641338 208266 641574
rect 208502 641338 208586 641574
rect 208822 641338 244266 641574
rect 244502 641338 244586 641574
rect 244822 641338 280266 641574
rect 280502 641338 280586 641574
rect 280822 641338 316266 641574
rect 316502 641338 316586 641574
rect 316822 641338 352266 641574
rect 352502 641338 352586 641574
rect 352822 641338 388266 641574
rect 388502 641338 388586 641574
rect 388822 641338 424266 641574
rect 424502 641338 424586 641574
rect 424822 641338 460266 641574
rect 460502 641338 460586 641574
rect 460822 641338 496266 641574
rect 496502 641338 496586 641574
rect 496822 641338 532266 641574
rect 532502 641338 532586 641574
rect 532822 641338 568266 641574
rect 568502 641338 568586 641574
rect 568822 641338 592062 641574
rect 592298 641338 592382 641574
rect 592618 641338 592650 641574
rect -8726 641306 592650 641338
rect -8726 638174 592650 638206
rect -8726 637938 -7734 638174
rect -7498 637938 -7414 638174
rect -7178 637938 24546 638174
rect 24782 637938 24866 638174
rect 25102 637938 60546 638174
rect 60782 637938 60866 638174
rect 61102 637938 96546 638174
rect 96782 637938 96866 638174
rect 97102 637938 132546 638174
rect 132782 637938 132866 638174
rect 133102 637938 168546 638174
rect 168782 637938 168866 638174
rect 169102 637938 204546 638174
rect 204782 637938 204866 638174
rect 205102 637938 240546 638174
rect 240782 637938 240866 638174
rect 241102 637938 276546 638174
rect 276782 637938 276866 638174
rect 277102 637938 312546 638174
rect 312782 637938 312866 638174
rect 313102 637938 348546 638174
rect 348782 637938 348866 638174
rect 349102 637938 384546 638174
rect 384782 637938 384866 638174
rect 385102 637938 420546 638174
rect 420782 637938 420866 638174
rect 421102 637938 456546 638174
rect 456782 637938 456866 638174
rect 457102 637938 492546 638174
rect 492782 637938 492866 638174
rect 493102 637938 528546 638174
rect 528782 637938 528866 638174
rect 529102 637938 564546 638174
rect 564782 637938 564866 638174
rect 565102 637938 591102 638174
rect 591338 637938 591422 638174
rect 591658 637938 592650 638174
rect -8726 637854 592650 637938
rect -8726 637618 -7734 637854
rect -7498 637618 -7414 637854
rect -7178 637618 24546 637854
rect 24782 637618 24866 637854
rect 25102 637618 60546 637854
rect 60782 637618 60866 637854
rect 61102 637618 96546 637854
rect 96782 637618 96866 637854
rect 97102 637618 132546 637854
rect 132782 637618 132866 637854
rect 133102 637618 168546 637854
rect 168782 637618 168866 637854
rect 169102 637618 204546 637854
rect 204782 637618 204866 637854
rect 205102 637618 240546 637854
rect 240782 637618 240866 637854
rect 241102 637618 276546 637854
rect 276782 637618 276866 637854
rect 277102 637618 312546 637854
rect 312782 637618 312866 637854
rect 313102 637618 348546 637854
rect 348782 637618 348866 637854
rect 349102 637618 384546 637854
rect 384782 637618 384866 637854
rect 385102 637618 420546 637854
rect 420782 637618 420866 637854
rect 421102 637618 456546 637854
rect 456782 637618 456866 637854
rect 457102 637618 492546 637854
rect 492782 637618 492866 637854
rect 493102 637618 528546 637854
rect 528782 637618 528866 637854
rect 529102 637618 564546 637854
rect 564782 637618 564866 637854
rect 565102 637618 591102 637854
rect 591338 637618 591422 637854
rect 591658 637618 592650 637854
rect -8726 637586 592650 637618
rect -8726 634454 592650 634486
rect -8726 634218 -6774 634454
rect -6538 634218 -6454 634454
rect -6218 634218 20826 634454
rect 21062 634218 21146 634454
rect 21382 634218 56826 634454
rect 57062 634218 57146 634454
rect 57382 634218 92826 634454
rect 93062 634218 93146 634454
rect 93382 634218 128826 634454
rect 129062 634218 129146 634454
rect 129382 634218 164826 634454
rect 165062 634218 165146 634454
rect 165382 634218 200826 634454
rect 201062 634218 201146 634454
rect 201382 634218 236826 634454
rect 237062 634218 237146 634454
rect 237382 634218 272826 634454
rect 273062 634218 273146 634454
rect 273382 634218 308826 634454
rect 309062 634218 309146 634454
rect 309382 634218 344826 634454
rect 345062 634218 345146 634454
rect 345382 634218 380826 634454
rect 381062 634218 381146 634454
rect 381382 634218 416826 634454
rect 417062 634218 417146 634454
rect 417382 634218 452826 634454
rect 453062 634218 453146 634454
rect 453382 634218 488826 634454
rect 489062 634218 489146 634454
rect 489382 634218 524826 634454
rect 525062 634218 525146 634454
rect 525382 634218 560826 634454
rect 561062 634218 561146 634454
rect 561382 634218 590142 634454
rect 590378 634218 590462 634454
rect 590698 634218 592650 634454
rect -8726 634134 592650 634218
rect -8726 633898 -6774 634134
rect -6538 633898 -6454 634134
rect -6218 633898 20826 634134
rect 21062 633898 21146 634134
rect 21382 633898 56826 634134
rect 57062 633898 57146 634134
rect 57382 633898 92826 634134
rect 93062 633898 93146 634134
rect 93382 633898 128826 634134
rect 129062 633898 129146 634134
rect 129382 633898 164826 634134
rect 165062 633898 165146 634134
rect 165382 633898 200826 634134
rect 201062 633898 201146 634134
rect 201382 633898 236826 634134
rect 237062 633898 237146 634134
rect 237382 633898 272826 634134
rect 273062 633898 273146 634134
rect 273382 633898 308826 634134
rect 309062 633898 309146 634134
rect 309382 633898 344826 634134
rect 345062 633898 345146 634134
rect 345382 633898 380826 634134
rect 381062 633898 381146 634134
rect 381382 633898 416826 634134
rect 417062 633898 417146 634134
rect 417382 633898 452826 634134
rect 453062 633898 453146 634134
rect 453382 633898 488826 634134
rect 489062 633898 489146 634134
rect 489382 633898 524826 634134
rect 525062 633898 525146 634134
rect 525382 633898 560826 634134
rect 561062 633898 561146 634134
rect 561382 633898 590142 634134
rect 590378 633898 590462 634134
rect 590698 633898 592650 634134
rect -8726 633866 592650 633898
rect -8726 630734 592650 630766
rect -8726 630498 -5814 630734
rect -5578 630498 -5494 630734
rect -5258 630498 17106 630734
rect 17342 630498 17426 630734
rect 17662 630498 53106 630734
rect 53342 630498 53426 630734
rect 53662 630498 89106 630734
rect 89342 630498 89426 630734
rect 89662 630498 125106 630734
rect 125342 630498 125426 630734
rect 125662 630498 161106 630734
rect 161342 630498 161426 630734
rect 161662 630498 197106 630734
rect 197342 630498 197426 630734
rect 197662 630498 233106 630734
rect 233342 630498 233426 630734
rect 233662 630498 269106 630734
rect 269342 630498 269426 630734
rect 269662 630498 305106 630734
rect 305342 630498 305426 630734
rect 305662 630498 341106 630734
rect 341342 630498 341426 630734
rect 341662 630498 377106 630734
rect 377342 630498 377426 630734
rect 377662 630498 413106 630734
rect 413342 630498 413426 630734
rect 413662 630498 449106 630734
rect 449342 630498 449426 630734
rect 449662 630498 485106 630734
rect 485342 630498 485426 630734
rect 485662 630498 521106 630734
rect 521342 630498 521426 630734
rect 521662 630498 557106 630734
rect 557342 630498 557426 630734
rect 557662 630498 589182 630734
rect 589418 630498 589502 630734
rect 589738 630498 592650 630734
rect -8726 630414 592650 630498
rect -8726 630178 -5814 630414
rect -5578 630178 -5494 630414
rect -5258 630178 17106 630414
rect 17342 630178 17426 630414
rect 17662 630178 53106 630414
rect 53342 630178 53426 630414
rect 53662 630178 89106 630414
rect 89342 630178 89426 630414
rect 89662 630178 125106 630414
rect 125342 630178 125426 630414
rect 125662 630178 161106 630414
rect 161342 630178 161426 630414
rect 161662 630178 197106 630414
rect 197342 630178 197426 630414
rect 197662 630178 233106 630414
rect 233342 630178 233426 630414
rect 233662 630178 269106 630414
rect 269342 630178 269426 630414
rect 269662 630178 305106 630414
rect 305342 630178 305426 630414
rect 305662 630178 341106 630414
rect 341342 630178 341426 630414
rect 341662 630178 377106 630414
rect 377342 630178 377426 630414
rect 377662 630178 413106 630414
rect 413342 630178 413426 630414
rect 413662 630178 449106 630414
rect 449342 630178 449426 630414
rect 449662 630178 485106 630414
rect 485342 630178 485426 630414
rect 485662 630178 521106 630414
rect 521342 630178 521426 630414
rect 521662 630178 557106 630414
rect 557342 630178 557426 630414
rect 557662 630178 589182 630414
rect 589418 630178 589502 630414
rect 589738 630178 592650 630414
rect -8726 630146 592650 630178
rect -8726 627014 592650 627046
rect -8726 626778 -4854 627014
rect -4618 626778 -4534 627014
rect -4298 626778 13386 627014
rect 13622 626778 13706 627014
rect 13942 626778 49386 627014
rect 49622 626778 49706 627014
rect 49942 626778 85386 627014
rect 85622 626778 85706 627014
rect 85942 626778 121386 627014
rect 121622 626778 121706 627014
rect 121942 626778 157386 627014
rect 157622 626778 157706 627014
rect 157942 626778 193386 627014
rect 193622 626778 193706 627014
rect 193942 626778 229386 627014
rect 229622 626778 229706 627014
rect 229942 626778 265386 627014
rect 265622 626778 265706 627014
rect 265942 626778 301386 627014
rect 301622 626778 301706 627014
rect 301942 626778 337386 627014
rect 337622 626778 337706 627014
rect 337942 626778 373386 627014
rect 373622 626778 373706 627014
rect 373942 626778 409386 627014
rect 409622 626778 409706 627014
rect 409942 626778 445386 627014
rect 445622 626778 445706 627014
rect 445942 626778 481386 627014
rect 481622 626778 481706 627014
rect 481942 626778 517386 627014
rect 517622 626778 517706 627014
rect 517942 626778 553386 627014
rect 553622 626778 553706 627014
rect 553942 626778 588222 627014
rect 588458 626778 588542 627014
rect 588778 626778 592650 627014
rect -8726 626694 592650 626778
rect -8726 626458 -4854 626694
rect -4618 626458 -4534 626694
rect -4298 626458 13386 626694
rect 13622 626458 13706 626694
rect 13942 626458 49386 626694
rect 49622 626458 49706 626694
rect 49942 626458 85386 626694
rect 85622 626458 85706 626694
rect 85942 626458 121386 626694
rect 121622 626458 121706 626694
rect 121942 626458 157386 626694
rect 157622 626458 157706 626694
rect 157942 626458 193386 626694
rect 193622 626458 193706 626694
rect 193942 626458 229386 626694
rect 229622 626458 229706 626694
rect 229942 626458 265386 626694
rect 265622 626458 265706 626694
rect 265942 626458 301386 626694
rect 301622 626458 301706 626694
rect 301942 626458 337386 626694
rect 337622 626458 337706 626694
rect 337942 626458 373386 626694
rect 373622 626458 373706 626694
rect 373942 626458 409386 626694
rect 409622 626458 409706 626694
rect 409942 626458 445386 626694
rect 445622 626458 445706 626694
rect 445942 626458 481386 626694
rect 481622 626458 481706 626694
rect 481942 626458 517386 626694
rect 517622 626458 517706 626694
rect 517942 626458 553386 626694
rect 553622 626458 553706 626694
rect 553942 626458 588222 626694
rect 588458 626458 588542 626694
rect 588778 626458 592650 626694
rect -8726 626426 592650 626458
rect -8726 623294 592650 623326
rect -8726 623058 -3894 623294
rect -3658 623058 -3574 623294
rect -3338 623058 9666 623294
rect 9902 623058 9986 623294
rect 10222 623058 45666 623294
rect 45902 623058 45986 623294
rect 46222 623058 81666 623294
rect 81902 623058 81986 623294
rect 82222 623058 117666 623294
rect 117902 623058 117986 623294
rect 118222 623058 153666 623294
rect 153902 623058 153986 623294
rect 154222 623058 189666 623294
rect 189902 623058 189986 623294
rect 190222 623058 225666 623294
rect 225902 623058 225986 623294
rect 226222 623058 261666 623294
rect 261902 623058 261986 623294
rect 262222 623058 297666 623294
rect 297902 623058 297986 623294
rect 298222 623058 333666 623294
rect 333902 623058 333986 623294
rect 334222 623058 369666 623294
rect 369902 623058 369986 623294
rect 370222 623058 405666 623294
rect 405902 623058 405986 623294
rect 406222 623058 441666 623294
rect 441902 623058 441986 623294
rect 442222 623058 477666 623294
rect 477902 623058 477986 623294
rect 478222 623058 513666 623294
rect 513902 623058 513986 623294
rect 514222 623058 549666 623294
rect 549902 623058 549986 623294
rect 550222 623058 587262 623294
rect 587498 623058 587582 623294
rect 587818 623058 592650 623294
rect -8726 622974 592650 623058
rect -8726 622738 -3894 622974
rect -3658 622738 -3574 622974
rect -3338 622738 9666 622974
rect 9902 622738 9986 622974
rect 10222 622738 45666 622974
rect 45902 622738 45986 622974
rect 46222 622738 81666 622974
rect 81902 622738 81986 622974
rect 82222 622738 117666 622974
rect 117902 622738 117986 622974
rect 118222 622738 153666 622974
rect 153902 622738 153986 622974
rect 154222 622738 189666 622974
rect 189902 622738 189986 622974
rect 190222 622738 225666 622974
rect 225902 622738 225986 622974
rect 226222 622738 261666 622974
rect 261902 622738 261986 622974
rect 262222 622738 297666 622974
rect 297902 622738 297986 622974
rect 298222 622738 333666 622974
rect 333902 622738 333986 622974
rect 334222 622738 369666 622974
rect 369902 622738 369986 622974
rect 370222 622738 405666 622974
rect 405902 622738 405986 622974
rect 406222 622738 441666 622974
rect 441902 622738 441986 622974
rect 442222 622738 477666 622974
rect 477902 622738 477986 622974
rect 478222 622738 513666 622974
rect 513902 622738 513986 622974
rect 514222 622738 549666 622974
rect 549902 622738 549986 622974
rect 550222 622738 587262 622974
rect 587498 622738 587582 622974
rect 587818 622738 592650 622974
rect -8726 622706 592650 622738
rect -8726 619574 592650 619606
rect -8726 619338 -2934 619574
rect -2698 619338 -2614 619574
rect -2378 619338 5946 619574
rect 6182 619338 6266 619574
rect 6502 619338 41946 619574
rect 42182 619338 42266 619574
rect 42502 619338 77946 619574
rect 78182 619338 78266 619574
rect 78502 619338 113946 619574
rect 114182 619338 114266 619574
rect 114502 619338 149946 619574
rect 150182 619338 150266 619574
rect 150502 619338 185946 619574
rect 186182 619338 186266 619574
rect 186502 619338 221946 619574
rect 222182 619338 222266 619574
rect 222502 619338 257946 619574
rect 258182 619338 258266 619574
rect 258502 619338 293946 619574
rect 294182 619338 294266 619574
rect 294502 619338 329946 619574
rect 330182 619338 330266 619574
rect 330502 619338 365946 619574
rect 366182 619338 366266 619574
rect 366502 619338 401946 619574
rect 402182 619338 402266 619574
rect 402502 619338 437946 619574
rect 438182 619338 438266 619574
rect 438502 619338 473946 619574
rect 474182 619338 474266 619574
rect 474502 619338 509946 619574
rect 510182 619338 510266 619574
rect 510502 619338 545946 619574
rect 546182 619338 546266 619574
rect 546502 619338 581946 619574
rect 582182 619338 582266 619574
rect 582502 619338 586302 619574
rect 586538 619338 586622 619574
rect 586858 619338 592650 619574
rect -8726 619254 592650 619338
rect -8726 619018 -2934 619254
rect -2698 619018 -2614 619254
rect -2378 619018 5946 619254
rect 6182 619018 6266 619254
rect 6502 619018 41946 619254
rect 42182 619018 42266 619254
rect 42502 619018 77946 619254
rect 78182 619018 78266 619254
rect 78502 619018 113946 619254
rect 114182 619018 114266 619254
rect 114502 619018 149946 619254
rect 150182 619018 150266 619254
rect 150502 619018 185946 619254
rect 186182 619018 186266 619254
rect 186502 619018 221946 619254
rect 222182 619018 222266 619254
rect 222502 619018 257946 619254
rect 258182 619018 258266 619254
rect 258502 619018 293946 619254
rect 294182 619018 294266 619254
rect 294502 619018 329946 619254
rect 330182 619018 330266 619254
rect 330502 619018 365946 619254
rect 366182 619018 366266 619254
rect 366502 619018 401946 619254
rect 402182 619018 402266 619254
rect 402502 619018 437946 619254
rect 438182 619018 438266 619254
rect 438502 619018 473946 619254
rect 474182 619018 474266 619254
rect 474502 619018 509946 619254
rect 510182 619018 510266 619254
rect 510502 619018 545946 619254
rect 546182 619018 546266 619254
rect 546502 619018 581946 619254
rect 582182 619018 582266 619254
rect 582502 619018 586302 619254
rect 586538 619018 586622 619254
rect 586858 619018 592650 619254
rect -8726 618986 592650 619018
rect -8726 615854 592650 615886
rect -8726 615618 -1974 615854
rect -1738 615618 -1654 615854
rect -1418 615618 2226 615854
rect 2462 615618 2546 615854
rect 2782 615618 38226 615854
rect 38462 615618 38546 615854
rect 38782 615618 74226 615854
rect 74462 615618 74546 615854
rect 74782 615618 110226 615854
rect 110462 615618 110546 615854
rect 110782 615618 146226 615854
rect 146462 615618 146546 615854
rect 146782 615618 182226 615854
rect 182462 615618 182546 615854
rect 182782 615618 218226 615854
rect 218462 615618 218546 615854
rect 218782 615618 254226 615854
rect 254462 615618 254546 615854
rect 254782 615618 290226 615854
rect 290462 615618 290546 615854
rect 290782 615618 326226 615854
rect 326462 615618 326546 615854
rect 326782 615618 362226 615854
rect 362462 615618 362546 615854
rect 362782 615618 398226 615854
rect 398462 615618 398546 615854
rect 398782 615618 434226 615854
rect 434462 615618 434546 615854
rect 434782 615618 470226 615854
rect 470462 615618 470546 615854
rect 470782 615618 506226 615854
rect 506462 615618 506546 615854
rect 506782 615618 542226 615854
rect 542462 615618 542546 615854
rect 542782 615618 578226 615854
rect 578462 615618 578546 615854
rect 578782 615618 585342 615854
rect 585578 615618 585662 615854
rect 585898 615618 592650 615854
rect -8726 615534 592650 615618
rect -8726 615298 -1974 615534
rect -1738 615298 -1654 615534
rect -1418 615298 2226 615534
rect 2462 615298 2546 615534
rect 2782 615298 38226 615534
rect 38462 615298 38546 615534
rect 38782 615298 74226 615534
rect 74462 615298 74546 615534
rect 74782 615298 110226 615534
rect 110462 615298 110546 615534
rect 110782 615298 146226 615534
rect 146462 615298 146546 615534
rect 146782 615298 182226 615534
rect 182462 615298 182546 615534
rect 182782 615298 218226 615534
rect 218462 615298 218546 615534
rect 218782 615298 254226 615534
rect 254462 615298 254546 615534
rect 254782 615298 290226 615534
rect 290462 615298 290546 615534
rect 290782 615298 326226 615534
rect 326462 615298 326546 615534
rect 326782 615298 362226 615534
rect 362462 615298 362546 615534
rect 362782 615298 398226 615534
rect 398462 615298 398546 615534
rect 398782 615298 434226 615534
rect 434462 615298 434546 615534
rect 434782 615298 470226 615534
rect 470462 615298 470546 615534
rect 470782 615298 506226 615534
rect 506462 615298 506546 615534
rect 506782 615298 542226 615534
rect 542462 615298 542546 615534
rect 542782 615298 578226 615534
rect 578462 615298 578546 615534
rect 578782 615298 585342 615534
rect 585578 615298 585662 615534
rect 585898 615298 592650 615534
rect -8726 615266 592650 615298
rect -8726 605894 592650 605926
rect -8726 605658 -8694 605894
rect -8458 605658 -8374 605894
rect -8138 605658 28266 605894
rect 28502 605658 28586 605894
rect 28822 605658 64266 605894
rect 64502 605658 64586 605894
rect 64822 605658 100266 605894
rect 100502 605658 100586 605894
rect 100822 605658 136266 605894
rect 136502 605658 136586 605894
rect 136822 605658 172266 605894
rect 172502 605658 172586 605894
rect 172822 605658 208266 605894
rect 208502 605658 208586 605894
rect 208822 605658 244266 605894
rect 244502 605658 244586 605894
rect 244822 605658 280266 605894
rect 280502 605658 280586 605894
rect 280822 605658 316266 605894
rect 316502 605658 316586 605894
rect 316822 605658 352266 605894
rect 352502 605658 352586 605894
rect 352822 605658 388266 605894
rect 388502 605658 388586 605894
rect 388822 605658 424266 605894
rect 424502 605658 424586 605894
rect 424822 605658 460266 605894
rect 460502 605658 460586 605894
rect 460822 605658 496266 605894
rect 496502 605658 496586 605894
rect 496822 605658 532266 605894
rect 532502 605658 532586 605894
rect 532822 605658 568266 605894
rect 568502 605658 568586 605894
rect 568822 605658 592062 605894
rect 592298 605658 592382 605894
rect 592618 605658 592650 605894
rect -8726 605574 592650 605658
rect -8726 605338 -8694 605574
rect -8458 605338 -8374 605574
rect -8138 605338 28266 605574
rect 28502 605338 28586 605574
rect 28822 605338 64266 605574
rect 64502 605338 64586 605574
rect 64822 605338 100266 605574
rect 100502 605338 100586 605574
rect 100822 605338 136266 605574
rect 136502 605338 136586 605574
rect 136822 605338 172266 605574
rect 172502 605338 172586 605574
rect 172822 605338 208266 605574
rect 208502 605338 208586 605574
rect 208822 605338 244266 605574
rect 244502 605338 244586 605574
rect 244822 605338 280266 605574
rect 280502 605338 280586 605574
rect 280822 605338 316266 605574
rect 316502 605338 316586 605574
rect 316822 605338 352266 605574
rect 352502 605338 352586 605574
rect 352822 605338 388266 605574
rect 388502 605338 388586 605574
rect 388822 605338 424266 605574
rect 424502 605338 424586 605574
rect 424822 605338 460266 605574
rect 460502 605338 460586 605574
rect 460822 605338 496266 605574
rect 496502 605338 496586 605574
rect 496822 605338 532266 605574
rect 532502 605338 532586 605574
rect 532822 605338 568266 605574
rect 568502 605338 568586 605574
rect 568822 605338 592062 605574
rect 592298 605338 592382 605574
rect 592618 605338 592650 605574
rect -8726 605306 592650 605338
rect -8726 602174 592650 602206
rect -8726 601938 -7734 602174
rect -7498 601938 -7414 602174
rect -7178 601938 24546 602174
rect 24782 601938 24866 602174
rect 25102 601938 60546 602174
rect 60782 601938 60866 602174
rect 61102 601938 96546 602174
rect 96782 601938 96866 602174
rect 97102 601938 132546 602174
rect 132782 601938 132866 602174
rect 133102 601938 168546 602174
rect 168782 601938 168866 602174
rect 169102 601938 204546 602174
rect 204782 601938 204866 602174
rect 205102 601938 240546 602174
rect 240782 601938 240866 602174
rect 241102 601938 276546 602174
rect 276782 601938 276866 602174
rect 277102 601938 312546 602174
rect 312782 601938 312866 602174
rect 313102 601938 348546 602174
rect 348782 601938 348866 602174
rect 349102 601938 384546 602174
rect 384782 601938 384866 602174
rect 385102 601938 420546 602174
rect 420782 601938 420866 602174
rect 421102 601938 456546 602174
rect 456782 601938 456866 602174
rect 457102 601938 492546 602174
rect 492782 601938 492866 602174
rect 493102 601938 528546 602174
rect 528782 601938 528866 602174
rect 529102 601938 564546 602174
rect 564782 601938 564866 602174
rect 565102 601938 591102 602174
rect 591338 601938 591422 602174
rect 591658 601938 592650 602174
rect -8726 601854 592650 601938
rect -8726 601618 -7734 601854
rect -7498 601618 -7414 601854
rect -7178 601618 24546 601854
rect 24782 601618 24866 601854
rect 25102 601618 60546 601854
rect 60782 601618 60866 601854
rect 61102 601618 96546 601854
rect 96782 601618 96866 601854
rect 97102 601618 132546 601854
rect 132782 601618 132866 601854
rect 133102 601618 168546 601854
rect 168782 601618 168866 601854
rect 169102 601618 204546 601854
rect 204782 601618 204866 601854
rect 205102 601618 240546 601854
rect 240782 601618 240866 601854
rect 241102 601618 276546 601854
rect 276782 601618 276866 601854
rect 277102 601618 312546 601854
rect 312782 601618 312866 601854
rect 313102 601618 348546 601854
rect 348782 601618 348866 601854
rect 349102 601618 384546 601854
rect 384782 601618 384866 601854
rect 385102 601618 420546 601854
rect 420782 601618 420866 601854
rect 421102 601618 456546 601854
rect 456782 601618 456866 601854
rect 457102 601618 492546 601854
rect 492782 601618 492866 601854
rect 493102 601618 528546 601854
rect 528782 601618 528866 601854
rect 529102 601618 564546 601854
rect 564782 601618 564866 601854
rect 565102 601618 591102 601854
rect 591338 601618 591422 601854
rect 591658 601618 592650 601854
rect -8726 601586 592650 601618
rect -8726 598454 592650 598486
rect -8726 598218 -6774 598454
rect -6538 598218 -6454 598454
rect -6218 598218 20826 598454
rect 21062 598218 21146 598454
rect 21382 598218 56826 598454
rect 57062 598218 57146 598454
rect 57382 598218 92826 598454
rect 93062 598218 93146 598454
rect 93382 598218 128826 598454
rect 129062 598218 129146 598454
rect 129382 598218 164826 598454
rect 165062 598218 165146 598454
rect 165382 598218 200826 598454
rect 201062 598218 201146 598454
rect 201382 598218 236826 598454
rect 237062 598218 237146 598454
rect 237382 598218 272826 598454
rect 273062 598218 273146 598454
rect 273382 598218 308826 598454
rect 309062 598218 309146 598454
rect 309382 598218 344826 598454
rect 345062 598218 345146 598454
rect 345382 598218 380826 598454
rect 381062 598218 381146 598454
rect 381382 598218 416826 598454
rect 417062 598218 417146 598454
rect 417382 598218 452826 598454
rect 453062 598218 453146 598454
rect 453382 598218 488826 598454
rect 489062 598218 489146 598454
rect 489382 598218 524826 598454
rect 525062 598218 525146 598454
rect 525382 598218 560826 598454
rect 561062 598218 561146 598454
rect 561382 598218 590142 598454
rect 590378 598218 590462 598454
rect 590698 598218 592650 598454
rect -8726 598134 592650 598218
rect -8726 597898 -6774 598134
rect -6538 597898 -6454 598134
rect -6218 597898 20826 598134
rect 21062 597898 21146 598134
rect 21382 597898 56826 598134
rect 57062 597898 57146 598134
rect 57382 597898 92826 598134
rect 93062 597898 93146 598134
rect 93382 597898 128826 598134
rect 129062 597898 129146 598134
rect 129382 597898 164826 598134
rect 165062 597898 165146 598134
rect 165382 597898 200826 598134
rect 201062 597898 201146 598134
rect 201382 597898 236826 598134
rect 237062 597898 237146 598134
rect 237382 597898 272826 598134
rect 273062 597898 273146 598134
rect 273382 597898 308826 598134
rect 309062 597898 309146 598134
rect 309382 597898 344826 598134
rect 345062 597898 345146 598134
rect 345382 597898 380826 598134
rect 381062 597898 381146 598134
rect 381382 597898 416826 598134
rect 417062 597898 417146 598134
rect 417382 597898 452826 598134
rect 453062 597898 453146 598134
rect 453382 597898 488826 598134
rect 489062 597898 489146 598134
rect 489382 597898 524826 598134
rect 525062 597898 525146 598134
rect 525382 597898 560826 598134
rect 561062 597898 561146 598134
rect 561382 597898 590142 598134
rect 590378 597898 590462 598134
rect 590698 597898 592650 598134
rect -8726 597866 592650 597898
rect -8726 594734 592650 594766
rect -8726 594498 -5814 594734
rect -5578 594498 -5494 594734
rect -5258 594498 17106 594734
rect 17342 594498 17426 594734
rect 17662 594498 53106 594734
rect 53342 594498 53426 594734
rect 53662 594498 89106 594734
rect 89342 594498 89426 594734
rect 89662 594498 125106 594734
rect 125342 594498 125426 594734
rect 125662 594498 161106 594734
rect 161342 594498 161426 594734
rect 161662 594498 197106 594734
rect 197342 594498 197426 594734
rect 197662 594498 233106 594734
rect 233342 594498 233426 594734
rect 233662 594498 269106 594734
rect 269342 594498 269426 594734
rect 269662 594498 305106 594734
rect 305342 594498 305426 594734
rect 305662 594498 341106 594734
rect 341342 594498 341426 594734
rect 341662 594498 377106 594734
rect 377342 594498 377426 594734
rect 377662 594498 413106 594734
rect 413342 594498 413426 594734
rect 413662 594498 449106 594734
rect 449342 594498 449426 594734
rect 449662 594498 485106 594734
rect 485342 594498 485426 594734
rect 485662 594498 521106 594734
rect 521342 594498 521426 594734
rect 521662 594498 557106 594734
rect 557342 594498 557426 594734
rect 557662 594498 589182 594734
rect 589418 594498 589502 594734
rect 589738 594498 592650 594734
rect -8726 594414 592650 594498
rect -8726 594178 -5814 594414
rect -5578 594178 -5494 594414
rect -5258 594178 17106 594414
rect 17342 594178 17426 594414
rect 17662 594178 53106 594414
rect 53342 594178 53426 594414
rect 53662 594178 89106 594414
rect 89342 594178 89426 594414
rect 89662 594178 125106 594414
rect 125342 594178 125426 594414
rect 125662 594178 161106 594414
rect 161342 594178 161426 594414
rect 161662 594178 197106 594414
rect 197342 594178 197426 594414
rect 197662 594178 233106 594414
rect 233342 594178 233426 594414
rect 233662 594178 269106 594414
rect 269342 594178 269426 594414
rect 269662 594178 305106 594414
rect 305342 594178 305426 594414
rect 305662 594178 341106 594414
rect 341342 594178 341426 594414
rect 341662 594178 377106 594414
rect 377342 594178 377426 594414
rect 377662 594178 413106 594414
rect 413342 594178 413426 594414
rect 413662 594178 449106 594414
rect 449342 594178 449426 594414
rect 449662 594178 485106 594414
rect 485342 594178 485426 594414
rect 485662 594178 521106 594414
rect 521342 594178 521426 594414
rect 521662 594178 557106 594414
rect 557342 594178 557426 594414
rect 557662 594178 589182 594414
rect 589418 594178 589502 594414
rect 589738 594178 592650 594414
rect -8726 594146 592650 594178
rect -8726 591014 592650 591046
rect -8726 590778 -4854 591014
rect -4618 590778 -4534 591014
rect -4298 590778 13386 591014
rect 13622 590778 13706 591014
rect 13942 590778 49386 591014
rect 49622 590778 49706 591014
rect 49942 590778 85386 591014
rect 85622 590778 85706 591014
rect 85942 590778 121386 591014
rect 121622 590778 121706 591014
rect 121942 590778 157386 591014
rect 157622 590778 157706 591014
rect 157942 590778 193386 591014
rect 193622 590778 193706 591014
rect 193942 590778 229386 591014
rect 229622 590778 229706 591014
rect 229942 590778 265386 591014
rect 265622 590778 265706 591014
rect 265942 590778 301386 591014
rect 301622 590778 301706 591014
rect 301942 590778 337386 591014
rect 337622 590778 337706 591014
rect 337942 590778 373386 591014
rect 373622 590778 373706 591014
rect 373942 590778 409386 591014
rect 409622 590778 409706 591014
rect 409942 590778 445386 591014
rect 445622 590778 445706 591014
rect 445942 590778 481386 591014
rect 481622 590778 481706 591014
rect 481942 590778 517386 591014
rect 517622 590778 517706 591014
rect 517942 590778 553386 591014
rect 553622 590778 553706 591014
rect 553942 590778 588222 591014
rect 588458 590778 588542 591014
rect 588778 590778 592650 591014
rect -8726 590694 592650 590778
rect -8726 590458 -4854 590694
rect -4618 590458 -4534 590694
rect -4298 590458 13386 590694
rect 13622 590458 13706 590694
rect 13942 590458 49386 590694
rect 49622 590458 49706 590694
rect 49942 590458 85386 590694
rect 85622 590458 85706 590694
rect 85942 590458 121386 590694
rect 121622 590458 121706 590694
rect 121942 590458 157386 590694
rect 157622 590458 157706 590694
rect 157942 590458 193386 590694
rect 193622 590458 193706 590694
rect 193942 590458 229386 590694
rect 229622 590458 229706 590694
rect 229942 590458 265386 590694
rect 265622 590458 265706 590694
rect 265942 590458 301386 590694
rect 301622 590458 301706 590694
rect 301942 590458 337386 590694
rect 337622 590458 337706 590694
rect 337942 590458 373386 590694
rect 373622 590458 373706 590694
rect 373942 590458 409386 590694
rect 409622 590458 409706 590694
rect 409942 590458 445386 590694
rect 445622 590458 445706 590694
rect 445942 590458 481386 590694
rect 481622 590458 481706 590694
rect 481942 590458 517386 590694
rect 517622 590458 517706 590694
rect 517942 590458 553386 590694
rect 553622 590458 553706 590694
rect 553942 590458 588222 590694
rect 588458 590458 588542 590694
rect 588778 590458 592650 590694
rect -8726 590426 592650 590458
rect -8726 587294 592650 587326
rect -8726 587058 -3894 587294
rect -3658 587058 -3574 587294
rect -3338 587058 9666 587294
rect 9902 587058 9986 587294
rect 10222 587058 45666 587294
rect 45902 587058 45986 587294
rect 46222 587058 81666 587294
rect 81902 587058 81986 587294
rect 82222 587058 117666 587294
rect 117902 587058 117986 587294
rect 118222 587058 153666 587294
rect 153902 587058 153986 587294
rect 154222 587058 189666 587294
rect 189902 587058 189986 587294
rect 190222 587058 225666 587294
rect 225902 587058 225986 587294
rect 226222 587058 261666 587294
rect 261902 587058 261986 587294
rect 262222 587058 297666 587294
rect 297902 587058 297986 587294
rect 298222 587058 333666 587294
rect 333902 587058 333986 587294
rect 334222 587058 369666 587294
rect 369902 587058 369986 587294
rect 370222 587058 405666 587294
rect 405902 587058 405986 587294
rect 406222 587058 441666 587294
rect 441902 587058 441986 587294
rect 442222 587058 477666 587294
rect 477902 587058 477986 587294
rect 478222 587058 513666 587294
rect 513902 587058 513986 587294
rect 514222 587058 549666 587294
rect 549902 587058 549986 587294
rect 550222 587058 587262 587294
rect 587498 587058 587582 587294
rect 587818 587058 592650 587294
rect -8726 586974 592650 587058
rect -8726 586738 -3894 586974
rect -3658 586738 -3574 586974
rect -3338 586738 9666 586974
rect 9902 586738 9986 586974
rect 10222 586738 45666 586974
rect 45902 586738 45986 586974
rect 46222 586738 81666 586974
rect 81902 586738 81986 586974
rect 82222 586738 117666 586974
rect 117902 586738 117986 586974
rect 118222 586738 153666 586974
rect 153902 586738 153986 586974
rect 154222 586738 189666 586974
rect 189902 586738 189986 586974
rect 190222 586738 225666 586974
rect 225902 586738 225986 586974
rect 226222 586738 261666 586974
rect 261902 586738 261986 586974
rect 262222 586738 297666 586974
rect 297902 586738 297986 586974
rect 298222 586738 333666 586974
rect 333902 586738 333986 586974
rect 334222 586738 369666 586974
rect 369902 586738 369986 586974
rect 370222 586738 405666 586974
rect 405902 586738 405986 586974
rect 406222 586738 441666 586974
rect 441902 586738 441986 586974
rect 442222 586738 477666 586974
rect 477902 586738 477986 586974
rect 478222 586738 513666 586974
rect 513902 586738 513986 586974
rect 514222 586738 549666 586974
rect 549902 586738 549986 586974
rect 550222 586738 587262 586974
rect 587498 586738 587582 586974
rect 587818 586738 592650 586974
rect -8726 586706 592650 586738
rect -8726 583574 592650 583606
rect -8726 583338 -2934 583574
rect -2698 583338 -2614 583574
rect -2378 583338 5946 583574
rect 6182 583338 6266 583574
rect 6502 583338 41946 583574
rect 42182 583338 42266 583574
rect 42502 583338 77946 583574
rect 78182 583338 78266 583574
rect 78502 583338 113946 583574
rect 114182 583338 114266 583574
rect 114502 583338 149946 583574
rect 150182 583338 150266 583574
rect 150502 583338 185946 583574
rect 186182 583338 186266 583574
rect 186502 583338 221946 583574
rect 222182 583338 222266 583574
rect 222502 583338 257946 583574
rect 258182 583338 258266 583574
rect 258502 583338 293946 583574
rect 294182 583338 294266 583574
rect 294502 583338 329946 583574
rect 330182 583338 330266 583574
rect 330502 583338 365946 583574
rect 366182 583338 366266 583574
rect 366502 583338 401946 583574
rect 402182 583338 402266 583574
rect 402502 583338 437946 583574
rect 438182 583338 438266 583574
rect 438502 583338 473946 583574
rect 474182 583338 474266 583574
rect 474502 583338 509946 583574
rect 510182 583338 510266 583574
rect 510502 583338 545946 583574
rect 546182 583338 546266 583574
rect 546502 583338 581946 583574
rect 582182 583338 582266 583574
rect 582502 583338 586302 583574
rect 586538 583338 586622 583574
rect 586858 583338 592650 583574
rect -8726 583254 592650 583338
rect -8726 583018 -2934 583254
rect -2698 583018 -2614 583254
rect -2378 583018 5946 583254
rect 6182 583018 6266 583254
rect 6502 583018 41946 583254
rect 42182 583018 42266 583254
rect 42502 583018 77946 583254
rect 78182 583018 78266 583254
rect 78502 583018 113946 583254
rect 114182 583018 114266 583254
rect 114502 583018 149946 583254
rect 150182 583018 150266 583254
rect 150502 583018 185946 583254
rect 186182 583018 186266 583254
rect 186502 583018 221946 583254
rect 222182 583018 222266 583254
rect 222502 583018 257946 583254
rect 258182 583018 258266 583254
rect 258502 583018 293946 583254
rect 294182 583018 294266 583254
rect 294502 583018 329946 583254
rect 330182 583018 330266 583254
rect 330502 583018 365946 583254
rect 366182 583018 366266 583254
rect 366502 583018 401946 583254
rect 402182 583018 402266 583254
rect 402502 583018 437946 583254
rect 438182 583018 438266 583254
rect 438502 583018 473946 583254
rect 474182 583018 474266 583254
rect 474502 583018 509946 583254
rect 510182 583018 510266 583254
rect 510502 583018 545946 583254
rect 546182 583018 546266 583254
rect 546502 583018 581946 583254
rect 582182 583018 582266 583254
rect 582502 583018 586302 583254
rect 586538 583018 586622 583254
rect 586858 583018 592650 583254
rect -8726 582986 592650 583018
rect -8726 579854 592650 579886
rect -8726 579618 -1974 579854
rect -1738 579618 -1654 579854
rect -1418 579618 2226 579854
rect 2462 579618 2546 579854
rect 2782 579618 38226 579854
rect 38462 579618 38546 579854
rect 38782 579618 74226 579854
rect 74462 579618 74546 579854
rect 74782 579618 110226 579854
rect 110462 579618 110546 579854
rect 110782 579618 146226 579854
rect 146462 579618 146546 579854
rect 146782 579618 182226 579854
rect 182462 579618 182546 579854
rect 182782 579618 218226 579854
rect 218462 579618 218546 579854
rect 218782 579618 254226 579854
rect 254462 579618 254546 579854
rect 254782 579618 290226 579854
rect 290462 579618 290546 579854
rect 290782 579618 326226 579854
rect 326462 579618 326546 579854
rect 326782 579618 362226 579854
rect 362462 579618 362546 579854
rect 362782 579618 398226 579854
rect 398462 579618 398546 579854
rect 398782 579618 434226 579854
rect 434462 579618 434546 579854
rect 434782 579618 470226 579854
rect 470462 579618 470546 579854
rect 470782 579618 506226 579854
rect 506462 579618 506546 579854
rect 506782 579618 542226 579854
rect 542462 579618 542546 579854
rect 542782 579618 578226 579854
rect 578462 579618 578546 579854
rect 578782 579618 585342 579854
rect 585578 579618 585662 579854
rect 585898 579618 592650 579854
rect -8726 579534 592650 579618
rect -8726 579298 -1974 579534
rect -1738 579298 -1654 579534
rect -1418 579298 2226 579534
rect 2462 579298 2546 579534
rect 2782 579298 38226 579534
rect 38462 579298 38546 579534
rect 38782 579298 74226 579534
rect 74462 579298 74546 579534
rect 74782 579298 110226 579534
rect 110462 579298 110546 579534
rect 110782 579298 146226 579534
rect 146462 579298 146546 579534
rect 146782 579298 182226 579534
rect 182462 579298 182546 579534
rect 182782 579298 218226 579534
rect 218462 579298 218546 579534
rect 218782 579298 254226 579534
rect 254462 579298 254546 579534
rect 254782 579298 290226 579534
rect 290462 579298 290546 579534
rect 290782 579298 326226 579534
rect 326462 579298 326546 579534
rect 326782 579298 362226 579534
rect 362462 579298 362546 579534
rect 362782 579298 398226 579534
rect 398462 579298 398546 579534
rect 398782 579298 434226 579534
rect 434462 579298 434546 579534
rect 434782 579298 470226 579534
rect 470462 579298 470546 579534
rect 470782 579298 506226 579534
rect 506462 579298 506546 579534
rect 506782 579298 542226 579534
rect 542462 579298 542546 579534
rect 542782 579298 578226 579534
rect 578462 579298 578546 579534
rect 578782 579298 585342 579534
rect 585578 579298 585662 579534
rect 585898 579298 592650 579534
rect -8726 579266 592650 579298
rect -8726 569894 592650 569926
rect -8726 569658 -8694 569894
rect -8458 569658 -8374 569894
rect -8138 569658 28266 569894
rect 28502 569658 28586 569894
rect 28822 569658 64266 569894
rect 64502 569658 64586 569894
rect 64822 569658 100266 569894
rect 100502 569658 100586 569894
rect 100822 569658 136266 569894
rect 136502 569658 136586 569894
rect 136822 569658 172266 569894
rect 172502 569658 172586 569894
rect 172822 569658 208266 569894
rect 208502 569658 208586 569894
rect 208822 569658 244266 569894
rect 244502 569658 244586 569894
rect 244822 569658 280266 569894
rect 280502 569658 280586 569894
rect 280822 569658 316266 569894
rect 316502 569658 316586 569894
rect 316822 569658 352266 569894
rect 352502 569658 352586 569894
rect 352822 569658 388266 569894
rect 388502 569658 388586 569894
rect 388822 569658 424266 569894
rect 424502 569658 424586 569894
rect 424822 569658 460266 569894
rect 460502 569658 460586 569894
rect 460822 569658 496266 569894
rect 496502 569658 496586 569894
rect 496822 569658 532266 569894
rect 532502 569658 532586 569894
rect 532822 569658 568266 569894
rect 568502 569658 568586 569894
rect 568822 569658 592062 569894
rect 592298 569658 592382 569894
rect 592618 569658 592650 569894
rect -8726 569574 592650 569658
rect -8726 569338 -8694 569574
rect -8458 569338 -8374 569574
rect -8138 569338 28266 569574
rect 28502 569338 28586 569574
rect 28822 569338 64266 569574
rect 64502 569338 64586 569574
rect 64822 569338 100266 569574
rect 100502 569338 100586 569574
rect 100822 569338 136266 569574
rect 136502 569338 136586 569574
rect 136822 569338 172266 569574
rect 172502 569338 172586 569574
rect 172822 569338 208266 569574
rect 208502 569338 208586 569574
rect 208822 569338 244266 569574
rect 244502 569338 244586 569574
rect 244822 569338 280266 569574
rect 280502 569338 280586 569574
rect 280822 569338 316266 569574
rect 316502 569338 316586 569574
rect 316822 569338 352266 569574
rect 352502 569338 352586 569574
rect 352822 569338 388266 569574
rect 388502 569338 388586 569574
rect 388822 569338 424266 569574
rect 424502 569338 424586 569574
rect 424822 569338 460266 569574
rect 460502 569338 460586 569574
rect 460822 569338 496266 569574
rect 496502 569338 496586 569574
rect 496822 569338 532266 569574
rect 532502 569338 532586 569574
rect 532822 569338 568266 569574
rect 568502 569338 568586 569574
rect 568822 569338 592062 569574
rect 592298 569338 592382 569574
rect 592618 569338 592650 569574
rect -8726 569306 592650 569338
rect -8726 566174 592650 566206
rect -8726 565938 -7734 566174
rect -7498 565938 -7414 566174
rect -7178 565938 24546 566174
rect 24782 565938 24866 566174
rect 25102 565938 60546 566174
rect 60782 565938 60866 566174
rect 61102 565938 96546 566174
rect 96782 565938 96866 566174
rect 97102 565938 132546 566174
rect 132782 565938 132866 566174
rect 133102 565938 168546 566174
rect 168782 565938 168866 566174
rect 169102 565938 204546 566174
rect 204782 565938 204866 566174
rect 205102 565938 240546 566174
rect 240782 565938 240866 566174
rect 241102 565938 276546 566174
rect 276782 565938 276866 566174
rect 277102 565938 312546 566174
rect 312782 565938 312866 566174
rect 313102 565938 348546 566174
rect 348782 565938 348866 566174
rect 349102 565938 384546 566174
rect 384782 565938 384866 566174
rect 385102 565938 420546 566174
rect 420782 565938 420866 566174
rect 421102 565938 456546 566174
rect 456782 565938 456866 566174
rect 457102 565938 492546 566174
rect 492782 565938 492866 566174
rect 493102 565938 528546 566174
rect 528782 565938 528866 566174
rect 529102 565938 564546 566174
rect 564782 565938 564866 566174
rect 565102 565938 591102 566174
rect 591338 565938 591422 566174
rect 591658 565938 592650 566174
rect -8726 565854 592650 565938
rect -8726 565618 -7734 565854
rect -7498 565618 -7414 565854
rect -7178 565618 24546 565854
rect 24782 565618 24866 565854
rect 25102 565618 60546 565854
rect 60782 565618 60866 565854
rect 61102 565618 96546 565854
rect 96782 565618 96866 565854
rect 97102 565618 132546 565854
rect 132782 565618 132866 565854
rect 133102 565618 168546 565854
rect 168782 565618 168866 565854
rect 169102 565618 204546 565854
rect 204782 565618 204866 565854
rect 205102 565618 240546 565854
rect 240782 565618 240866 565854
rect 241102 565618 276546 565854
rect 276782 565618 276866 565854
rect 277102 565618 312546 565854
rect 312782 565618 312866 565854
rect 313102 565618 348546 565854
rect 348782 565618 348866 565854
rect 349102 565618 384546 565854
rect 384782 565618 384866 565854
rect 385102 565618 420546 565854
rect 420782 565618 420866 565854
rect 421102 565618 456546 565854
rect 456782 565618 456866 565854
rect 457102 565618 492546 565854
rect 492782 565618 492866 565854
rect 493102 565618 528546 565854
rect 528782 565618 528866 565854
rect 529102 565618 564546 565854
rect 564782 565618 564866 565854
rect 565102 565618 591102 565854
rect 591338 565618 591422 565854
rect 591658 565618 592650 565854
rect -8726 565586 592650 565618
rect -8726 562454 592650 562486
rect -8726 562218 -6774 562454
rect -6538 562218 -6454 562454
rect -6218 562218 20826 562454
rect 21062 562218 21146 562454
rect 21382 562218 56826 562454
rect 57062 562218 57146 562454
rect 57382 562218 92826 562454
rect 93062 562218 93146 562454
rect 93382 562218 128826 562454
rect 129062 562218 129146 562454
rect 129382 562218 164826 562454
rect 165062 562218 165146 562454
rect 165382 562218 200826 562454
rect 201062 562218 201146 562454
rect 201382 562218 236826 562454
rect 237062 562218 237146 562454
rect 237382 562218 272826 562454
rect 273062 562218 273146 562454
rect 273382 562218 308826 562454
rect 309062 562218 309146 562454
rect 309382 562218 344826 562454
rect 345062 562218 345146 562454
rect 345382 562218 380826 562454
rect 381062 562218 381146 562454
rect 381382 562218 416826 562454
rect 417062 562218 417146 562454
rect 417382 562218 452826 562454
rect 453062 562218 453146 562454
rect 453382 562218 488826 562454
rect 489062 562218 489146 562454
rect 489382 562218 524826 562454
rect 525062 562218 525146 562454
rect 525382 562218 560826 562454
rect 561062 562218 561146 562454
rect 561382 562218 590142 562454
rect 590378 562218 590462 562454
rect 590698 562218 592650 562454
rect -8726 562134 592650 562218
rect -8726 561898 -6774 562134
rect -6538 561898 -6454 562134
rect -6218 561898 20826 562134
rect 21062 561898 21146 562134
rect 21382 561898 56826 562134
rect 57062 561898 57146 562134
rect 57382 561898 92826 562134
rect 93062 561898 93146 562134
rect 93382 561898 128826 562134
rect 129062 561898 129146 562134
rect 129382 561898 164826 562134
rect 165062 561898 165146 562134
rect 165382 561898 200826 562134
rect 201062 561898 201146 562134
rect 201382 561898 236826 562134
rect 237062 561898 237146 562134
rect 237382 561898 272826 562134
rect 273062 561898 273146 562134
rect 273382 561898 308826 562134
rect 309062 561898 309146 562134
rect 309382 561898 344826 562134
rect 345062 561898 345146 562134
rect 345382 561898 380826 562134
rect 381062 561898 381146 562134
rect 381382 561898 416826 562134
rect 417062 561898 417146 562134
rect 417382 561898 452826 562134
rect 453062 561898 453146 562134
rect 453382 561898 488826 562134
rect 489062 561898 489146 562134
rect 489382 561898 524826 562134
rect 525062 561898 525146 562134
rect 525382 561898 560826 562134
rect 561062 561898 561146 562134
rect 561382 561898 590142 562134
rect 590378 561898 590462 562134
rect 590698 561898 592650 562134
rect -8726 561866 592650 561898
rect -8726 558734 592650 558766
rect -8726 558498 -5814 558734
rect -5578 558498 -5494 558734
rect -5258 558498 17106 558734
rect 17342 558498 17426 558734
rect 17662 558498 53106 558734
rect 53342 558498 53426 558734
rect 53662 558498 89106 558734
rect 89342 558498 89426 558734
rect 89662 558498 125106 558734
rect 125342 558498 125426 558734
rect 125662 558498 161106 558734
rect 161342 558498 161426 558734
rect 161662 558498 197106 558734
rect 197342 558498 197426 558734
rect 197662 558498 233106 558734
rect 233342 558498 233426 558734
rect 233662 558498 269106 558734
rect 269342 558498 269426 558734
rect 269662 558498 305106 558734
rect 305342 558498 305426 558734
rect 305662 558498 341106 558734
rect 341342 558498 341426 558734
rect 341662 558498 377106 558734
rect 377342 558498 377426 558734
rect 377662 558498 413106 558734
rect 413342 558498 413426 558734
rect 413662 558498 449106 558734
rect 449342 558498 449426 558734
rect 449662 558498 485106 558734
rect 485342 558498 485426 558734
rect 485662 558498 521106 558734
rect 521342 558498 521426 558734
rect 521662 558498 557106 558734
rect 557342 558498 557426 558734
rect 557662 558498 589182 558734
rect 589418 558498 589502 558734
rect 589738 558498 592650 558734
rect -8726 558414 592650 558498
rect -8726 558178 -5814 558414
rect -5578 558178 -5494 558414
rect -5258 558178 17106 558414
rect 17342 558178 17426 558414
rect 17662 558178 53106 558414
rect 53342 558178 53426 558414
rect 53662 558178 89106 558414
rect 89342 558178 89426 558414
rect 89662 558178 125106 558414
rect 125342 558178 125426 558414
rect 125662 558178 161106 558414
rect 161342 558178 161426 558414
rect 161662 558178 197106 558414
rect 197342 558178 197426 558414
rect 197662 558178 233106 558414
rect 233342 558178 233426 558414
rect 233662 558178 269106 558414
rect 269342 558178 269426 558414
rect 269662 558178 305106 558414
rect 305342 558178 305426 558414
rect 305662 558178 341106 558414
rect 341342 558178 341426 558414
rect 341662 558178 377106 558414
rect 377342 558178 377426 558414
rect 377662 558178 413106 558414
rect 413342 558178 413426 558414
rect 413662 558178 449106 558414
rect 449342 558178 449426 558414
rect 449662 558178 485106 558414
rect 485342 558178 485426 558414
rect 485662 558178 521106 558414
rect 521342 558178 521426 558414
rect 521662 558178 557106 558414
rect 557342 558178 557426 558414
rect 557662 558178 589182 558414
rect 589418 558178 589502 558414
rect 589738 558178 592650 558414
rect -8726 558146 592650 558178
rect -8726 555014 592650 555046
rect -8726 554778 -4854 555014
rect -4618 554778 -4534 555014
rect -4298 554778 13386 555014
rect 13622 554778 13706 555014
rect 13942 554778 49386 555014
rect 49622 554778 49706 555014
rect 49942 554778 85386 555014
rect 85622 554778 85706 555014
rect 85942 554778 121386 555014
rect 121622 554778 121706 555014
rect 121942 554778 157386 555014
rect 157622 554778 157706 555014
rect 157942 554778 193386 555014
rect 193622 554778 193706 555014
rect 193942 554778 229386 555014
rect 229622 554778 229706 555014
rect 229942 554778 265386 555014
rect 265622 554778 265706 555014
rect 265942 554778 301386 555014
rect 301622 554778 301706 555014
rect 301942 554778 337386 555014
rect 337622 554778 337706 555014
rect 337942 554778 373386 555014
rect 373622 554778 373706 555014
rect 373942 554778 409386 555014
rect 409622 554778 409706 555014
rect 409942 554778 445386 555014
rect 445622 554778 445706 555014
rect 445942 554778 481386 555014
rect 481622 554778 481706 555014
rect 481942 554778 517386 555014
rect 517622 554778 517706 555014
rect 517942 554778 553386 555014
rect 553622 554778 553706 555014
rect 553942 554778 588222 555014
rect 588458 554778 588542 555014
rect 588778 554778 592650 555014
rect -8726 554694 592650 554778
rect -8726 554458 -4854 554694
rect -4618 554458 -4534 554694
rect -4298 554458 13386 554694
rect 13622 554458 13706 554694
rect 13942 554458 49386 554694
rect 49622 554458 49706 554694
rect 49942 554458 85386 554694
rect 85622 554458 85706 554694
rect 85942 554458 121386 554694
rect 121622 554458 121706 554694
rect 121942 554458 157386 554694
rect 157622 554458 157706 554694
rect 157942 554458 193386 554694
rect 193622 554458 193706 554694
rect 193942 554458 229386 554694
rect 229622 554458 229706 554694
rect 229942 554458 265386 554694
rect 265622 554458 265706 554694
rect 265942 554458 301386 554694
rect 301622 554458 301706 554694
rect 301942 554458 337386 554694
rect 337622 554458 337706 554694
rect 337942 554458 373386 554694
rect 373622 554458 373706 554694
rect 373942 554458 409386 554694
rect 409622 554458 409706 554694
rect 409942 554458 445386 554694
rect 445622 554458 445706 554694
rect 445942 554458 481386 554694
rect 481622 554458 481706 554694
rect 481942 554458 517386 554694
rect 517622 554458 517706 554694
rect 517942 554458 553386 554694
rect 553622 554458 553706 554694
rect 553942 554458 588222 554694
rect 588458 554458 588542 554694
rect 588778 554458 592650 554694
rect -8726 554426 592650 554458
rect -8726 551294 592650 551326
rect -8726 551058 -3894 551294
rect -3658 551058 -3574 551294
rect -3338 551058 9666 551294
rect 9902 551058 9986 551294
rect 10222 551058 45666 551294
rect 45902 551058 45986 551294
rect 46222 551058 81666 551294
rect 81902 551058 81986 551294
rect 82222 551058 117666 551294
rect 117902 551058 117986 551294
rect 118222 551058 153666 551294
rect 153902 551058 153986 551294
rect 154222 551058 189666 551294
rect 189902 551058 189986 551294
rect 190222 551058 225666 551294
rect 225902 551058 225986 551294
rect 226222 551058 261666 551294
rect 261902 551058 261986 551294
rect 262222 551058 297666 551294
rect 297902 551058 297986 551294
rect 298222 551058 333666 551294
rect 333902 551058 333986 551294
rect 334222 551058 369666 551294
rect 369902 551058 369986 551294
rect 370222 551058 405666 551294
rect 405902 551058 405986 551294
rect 406222 551058 441666 551294
rect 441902 551058 441986 551294
rect 442222 551058 477666 551294
rect 477902 551058 477986 551294
rect 478222 551058 513666 551294
rect 513902 551058 513986 551294
rect 514222 551058 549666 551294
rect 549902 551058 549986 551294
rect 550222 551058 587262 551294
rect 587498 551058 587582 551294
rect 587818 551058 592650 551294
rect -8726 550974 592650 551058
rect -8726 550738 -3894 550974
rect -3658 550738 -3574 550974
rect -3338 550738 9666 550974
rect 9902 550738 9986 550974
rect 10222 550738 45666 550974
rect 45902 550738 45986 550974
rect 46222 550738 81666 550974
rect 81902 550738 81986 550974
rect 82222 550738 117666 550974
rect 117902 550738 117986 550974
rect 118222 550738 153666 550974
rect 153902 550738 153986 550974
rect 154222 550738 189666 550974
rect 189902 550738 189986 550974
rect 190222 550738 225666 550974
rect 225902 550738 225986 550974
rect 226222 550738 261666 550974
rect 261902 550738 261986 550974
rect 262222 550738 297666 550974
rect 297902 550738 297986 550974
rect 298222 550738 333666 550974
rect 333902 550738 333986 550974
rect 334222 550738 369666 550974
rect 369902 550738 369986 550974
rect 370222 550738 405666 550974
rect 405902 550738 405986 550974
rect 406222 550738 441666 550974
rect 441902 550738 441986 550974
rect 442222 550738 477666 550974
rect 477902 550738 477986 550974
rect 478222 550738 513666 550974
rect 513902 550738 513986 550974
rect 514222 550738 549666 550974
rect 549902 550738 549986 550974
rect 550222 550738 587262 550974
rect 587498 550738 587582 550974
rect 587818 550738 592650 550974
rect -8726 550706 592650 550738
rect -8726 547574 592650 547606
rect -8726 547338 -2934 547574
rect -2698 547338 -2614 547574
rect -2378 547338 5946 547574
rect 6182 547338 6266 547574
rect 6502 547338 41946 547574
rect 42182 547338 42266 547574
rect 42502 547338 77946 547574
rect 78182 547338 78266 547574
rect 78502 547338 113946 547574
rect 114182 547338 114266 547574
rect 114502 547338 149946 547574
rect 150182 547338 150266 547574
rect 150502 547338 185946 547574
rect 186182 547338 186266 547574
rect 186502 547338 221946 547574
rect 222182 547338 222266 547574
rect 222502 547338 257946 547574
rect 258182 547338 258266 547574
rect 258502 547338 293946 547574
rect 294182 547338 294266 547574
rect 294502 547338 329946 547574
rect 330182 547338 330266 547574
rect 330502 547338 365946 547574
rect 366182 547338 366266 547574
rect 366502 547338 401946 547574
rect 402182 547338 402266 547574
rect 402502 547338 437946 547574
rect 438182 547338 438266 547574
rect 438502 547338 473946 547574
rect 474182 547338 474266 547574
rect 474502 547338 509946 547574
rect 510182 547338 510266 547574
rect 510502 547338 545946 547574
rect 546182 547338 546266 547574
rect 546502 547338 581946 547574
rect 582182 547338 582266 547574
rect 582502 547338 586302 547574
rect 586538 547338 586622 547574
rect 586858 547338 592650 547574
rect -8726 547254 592650 547338
rect -8726 547018 -2934 547254
rect -2698 547018 -2614 547254
rect -2378 547018 5946 547254
rect 6182 547018 6266 547254
rect 6502 547018 41946 547254
rect 42182 547018 42266 547254
rect 42502 547018 77946 547254
rect 78182 547018 78266 547254
rect 78502 547018 113946 547254
rect 114182 547018 114266 547254
rect 114502 547018 149946 547254
rect 150182 547018 150266 547254
rect 150502 547018 185946 547254
rect 186182 547018 186266 547254
rect 186502 547018 221946 547254
rect 222182 547018 222266 547254
rect 222502 547018 257946 547254
rect 258182 547018 258266 547254
rect 258502 547018 293946 547254
rect 294182 547018 294266 547254
rect 294502 547018 329946 547254
rect 330182 547018 330266 547254
rect 330502 547018 365946 547254
rect 366182 547018 366266 547254
rect 366502 547018 401946 547254
rect 402182 547018 402266 547254
rect 402502 547018 437946 547254
rect 438182 547018 438266 547254
rect 438502 547018 473946 547254
rect 474182 547018 474266 547254
rect 474502 547018 509946 547254
rect 510182 547018 510266 547254
rect 510502 547018 545946 547254
rect 546182 547018 546266 547254
rect 546502 547018 581946 547254
rect 582182 547018 582266 547254
rect 582502 547018 586302 547254
rect 586538 547018 586622 547254
rect 586858 547018 592650 547254
rect -8726 546986 592650 547018
rect -8726 543854 592650 543886
rect -8726 543618 -1974 543854
rect -1738 543618 -1654 543854
rect -1418 543618 2226 543854
rect 2462 543618 2546 543854
rect 2782 543618 38226 543854
rect 38462 543618 38546 543854
rect 38782 543618 74226 543854
rect 74462 543618 74546 543854
rect 74782 543618 110226 543854
rect 110462 543618 110546 543854
rect 110782 543618 146226 543854
rect 146462 543618 146546 543854
rect 146782 543618 182226 543854
rect 182462 543618 182546 543854
rect 182782 543618 218226 543854
rect 218462 543618 218546 543854
rect 218782 543618 254226 543854
rect 254462 543618 254546 543854
rect 254782 543618 290226 543854
rect 290462 543618 290546 543854
rect 290782 543618 326226 543854
rect 326462 543618 326546 543854
rect 326782 543618 362226 543854
rect 362462 543618 362546 543854
rect 362782 543618 398226 543854
rect 398462 543618 398546 543854
rect 398782 543618 434226 543854
rect 434462 543618 434546 543854
rect 434782 543618 470226 543854
rect 470462 543618 470546 543854
rect 470782 543618 506226 543854
rect 506462 543618 506546 543854
rect 506782 543618 542226 543854
rect 542462 543618 542546 543854
rect 542782 543618 578226 543854
rect 578462 543618 578546 543854
rect 578782 543618 585342 543854
rect 585578 543618 585662 543854
rect 585898 543618 592650 543854
rect -8726 543534 592650 543618
rect -8726 543298 -1974 543534
rect -1738 543298 -1654 543534
rect -1418 543298 2226 543534
rect 2462 543298 2546 543534
rect 2782 543298 38226 543534
rect 38462 543298 38546 543534
rect 38782 543298 74226 543534
rect 74462 543298 74546 543534
rect 74782 543298 110226 543534
rect 110462 543298 110546 543534
rect 110782 543298 146226 543534
rect 146462 543298 146546 543534
rect 146782 543298 182226 543534
rect 182462 543298 182546 543534
rect 182782 543298 218226 543534
rect 218462 543298 218546 543534
rect 218782 543298 254226 543534
rect 254462 543298 254546 543534
rect 254782 543298 290226 543534
rect 290462 543298 290546 543534
rect 290782 543298 326226 543534
rect 326462 543298 326546 543534
rect 326782 543298 362226 543534
rect 362462 543298 362546 543534
rect 362782 543298 398226 543534
rect 398462 543298 398546 543534
rect 398782 543298 434226 543534
rect 434462 543298 434546 543534
rect 434782 543298 470226 543534
rect 470462 543298 470546 543534
rect 470782 543298 506226 543534
rect 506462 543298 506546 543534
rect 506782 543298 542226 543534
rect 542462 543298 542546 543534
rect 542782 543298 578226 543534
rect 578462 543298 578546 543534
rect 578782 543298 585342 543534
rect 585578 543298 585662 543534
rect 585898 543298 592650 543534
rect -8726 543266 592650 543298
rect -8726 533894 592650 533926
rect -8726 533658 -8694 533894
rect -8458 533658 -8374 533894
rect -8138 533658 28266 533894
rect 28502 533658 28586 533894
rect 28822 533658 64266 533894
rect 64502 533658 64586 533894
rect 64822 533658 100266 533894
rect 100502 533658 100586 533894
rect 100822 533658 136266 533894
rect 136502 533658 136586 533894
rect 136822 533658 172266 533894
rect 172502 533658 172586 533894
rect 172822 533658 208266 533894
rect 208502 533658 208586 533894
rect 208822 533658 244266 533894
rect 244502 533658 244586 533894
rect 244822 533658 280266 533894
rect 280502 533658 280586 533894
rect 280822 533658 316266 533894
rect 316502 533658 316586 533894
rect 316822 533658 352266 533894
rect 352502 533658 352586 533894
rect 352822 533658 388266 533894
rect 388502 533658 388586 533894
rect 388822 533658 424266 533894
rect 424502 533658 424586 533894
rect 424822 533658 460266 533894
rect 460502 533658 460586 533894
rect 460822 533658 496266 533894
rect 496502 533658 496586 533894
rect 496822 533658 532266 533894
rect 532502 533658 532586 533894
rect 532822 533658 568266 533894
rect 568502 533658 568586 533894
rect 568822 533658 592062 533894
rect 592298 533658 592382 533894
rect 592618 533658 592650 533894
rect -8726 533574 592650 533658
rect -8726 533338 -8694 533574
rect -8458 533338 -8374 533574
rect -8138 533338 28266 533574
rect 28502 533338 28586 533574
rect 28822 533338 64266 533574
rect 64502 533338 64586 533574
rect 64822 533338 100266 533574
rect 100502 533338 100586 533574
rect 100822 533338 136266 533574
rect 136502 533338 136586 533574
rect 136822 533338 172266 533574
rect 172502 533338 172586 533574
rect 172822 533338 208266 533574
rect 208502 533338 208586 533574
rect 208822 533338 244266 533574
rect 244502 533338 244586 533574
rect 244822 533338 280266 533574
rect 280502 533338 280586 533574
rect 280822 533338 316266 533574
rect 316502 533338 316586 533574
rect 316822 533338 352266 533574
rect 352502 533338 352586 533574
rect 352822 533338 388266 533574
rect 388502 533338 388586 533574
rect 388822 533338 424266 533574
rect 424502 533338 424586 533574
rect 424822 533338 460266 533574
rect 460502 533338 460586 533574
rect 460822 533338 496266 533574
rect 496502 533338 496586 533574
rect 496822 533338 532266 533574
rect 532502 533338 532586 533574
rect 532822 533338 568266 533574
rect 568502 533338 568586 533574
rect 568822 533338 592062 533574
rect 592298 533338 592382 533574
rect 592618 533338 592650 533574
rect -8726 533306 592650 533338
rect -8726 530174 592650 530206
rect -8726 529938 -7734 530174
rect -7498 529938 -7414 530174
rect -7178 529938 24546 530174
rect 24782 529938 24866 530174
rect 25102 529938 60546 530174
rect 60782 529938 60866 530174
rect 61102 529938 96546 530174
rect 96782 529938 96866 530174
rect 97102 529938 132546 530174
rect 132782 529938 132866 530174
rect 133102 529938 168546 530174
rect 168782 529938 168866 530174
rect 169102 529938 204546 530174
rect 204782 529938 204866 530174
rect 205102 529938 240546 530174
rect 240782 529938 240866 530174
rect 241102 529938 276546 530174
rect 276782 529938 276866 530174
rect 277102 529938 312546 530174
rect 312782 529938 312866 530174
rect 313102 529938 348546 530174
rect 348782 529938 348866 530174
rect 349102 529938 384546 530174
rect 384782 529938 384866 530174
rect 385102 529938 420546 530174
rect 420782 529938 420866 530174
rect 421102 529938 456546 530174
rect 456782 529938 456866 530174
rect 457102 529938 492546 530174
rect 492782 529938 492866 530174
rect 493102 529938 528546 530174
rect 528782 529938 528866 530174
rect 529102 529938 564546 530174
rect 564782 529938 564866 530174
rect 565102 529938 591102 530174
rect 591338 529938 591422 530174
rect 591658 529938 592650 530174
rect -8726 529854 592650 529938
rect -8726 529618 -7734 529854
rect -7498 529618 -7414 529854
rect -7178 529618 24546 529854
rect 24782 529618 24866 529854
rect 25102 529618 60546 529854
rect 60782 529618 60866 529854
rect 61102 529618 96546 529854
rect 96782 529618 96866 529854
rect 97102 529618 132546 529854
rect 132782 529618 132866 529854
rect 133102 529618 168546 529854
rect 168782 529618 168866 529854
rect 169102 529618 204546 529854
rect 204782 529618 204866 529854
rect 205102 529618 240546 529854
rect 240782 529618 240866 529854
rect 241102 529618 276546 529854
rect 276782 529618 276866 529854
rect 277102 529618 312546 529854
rect 312782 529618 312866 529854
rect 313102 529618 348546 529854
rect 348782 529618 348866 529854
rect 349102 529618 384546 529854
rect 384782 529618 384866 529854
rect 385102 529618 420546 529854
rect 420782 529618 420866 529854
rect 421102 529618 456546 529854
rect 456782 529618 456866 529854
rect 457102 529618 492546 529854
rect 492782 529618 492866 529854
rect 493102 529618 528546 529854
rect 528782 529618 528866 529854
rect 529102 529618 564546 529854
rect 564782 529618 564866 529854
rect 565102 529618 591102 529854
rect 591338 529618 591422 529854
rect 591658 529618 592650 529854
rect -8726 529586 592650 529618
rect -8726 526454 592650 526486
rect -8726 526218 -6774 526454
rect -6538 526218 -6454 526454
rect -6218 526218 20826 526454
rect 21062 526218 21146 526454
rect 21382 526218 56826 526454
rect 57062 526218 57146 526454
rect 57382 526218 92826 526454
rect 93062 526218 93146 526454
rect 93382 526218 128826 526454
rect 129062 526218 129146 526454
rect 129382 526218 164826 526454
rect 165062 526218 165146 526454
rect 165382 526218 200826 526454
rect 201062 526218 201146 526454
rect 201382 526218 236826 526454
rect 237062 526218 237146 526454
rect 237382 526218 272826 526454
rect 273062 526218 273146 526454
rect 273382 526218 308826 526454
rect 309062 526218 309146 526454
rect 309382 526218 344826 526454
rect 345062 526218 345146 526454
rect 345382 526218 380826 526454
rect 381062 526218 381146 526454
rect 381382 526218 416826 526454
rect 417062 526218 417146 526454
rect 417382 526218 452826 526454
rect 453062 526218 453146 526454
rect 453382 526218 488826 526454
rect 489062 526218 489146 526454
rect 489382 526218 524826 526454
rect 525062 526218 525146 526454
rect 525382 526218 560826 526454
rect 561062 526218 561146 526454
rect 561382 526218 590142 526454
rect 590378 526218 590462 526454
rect 590698 526218 592650 526454
rect -8726 526134 592650 526218
rect -8726 525898 -6774 526134
rect -6538 525898 -6454 526134
rect -6218 525898 20826 526134
rect 21062 525898 21146 526134
rect 21382 525898 56826 526134
rect 57062 525898 57146 526134
rect 57382 525898 92826 526134
rect 93062 525898 93146 526134
rect 93382 525898 128826 526134
rect 129062 525898 129146 526134
rect 129382 525898 164826 526134
rect 165062 525898 165146 526134
rect 165382 525898 200826 526134
rect 201062 525898 201146 526134
rect 201382 525898 236826 526134
rect 237062 525898 237146 526134
rect 237382 525898 272826 526134
rect 273062 525898 273146 526134
rect 273382 525898 308826 526134
rect 309062 525898 309146 526134
rect 309382 525898 344826 526134
rect 345062 525898 345146 526134
rect 345382 525898 380826 526134
rect 381062 525898 381146 526134
rect 381382 525898 416826 526134
rect 417062 525898 417146 526134
rect 417382 525898 452826 526134
rect 453062 525898 453146 526134
rect 453382 525898 488826 526134
rect 489062 525898 489146 526134
rect 489382 525898 524826 526134
rect 525062 525898 525146 526134
rect 525382 525898 560826 526134
rect 561062 525898 561146 526134
rect 561382 525898 590142 526134
rect 590378 525898 590462 526134
rect 590698 525898 592650 526134
rect -8726 525866 592650 525898
rect -8726 522734 592650 522766
rect -8726 522498 -5814 522734
rect -5578 522498 -5494 522734
rect -5258 522498 17106 522734
rect 17342 522498 17426 522734
rect 17662 522498 53106 522734
rect 53342 522498 53426 522734
rect 53662 522498 89106 522734
rect 89342 522498 89426 522734
rect 89662 522498 125106 522734
rect 125342 522498 125426 522734
rect 125662 522498 161106 522734
rect 161342 522498 161426 522734
rect 161662 522498 197106 522734
rect 197342 522498 197426 522734
rect 197662 522498 233106 522734
rect 233342 522498 233426 522734
rect 233662 522498 269106 522734
rect 269342 522498 269426 522734
rect 269662 522498 305106 522734
rect 305342 522498 305426 522734
rect 305662 522498 341106 522734
rect 341342 522498 341426 522734
rect 341662 522498 377106 522734
rect 377342 522498 377426 522734
rect 377662 522498 413106 522734
rect 413342 522498 413426 522734
rect 413662 522498 449106 522734
rect 449342 522498 449426 522734
rect 449662 522498 485106 522734
rect 485342 522498 485426 522734
rect 485662 522498 521106 522734
rect 521342 522498 521426 522734
rect 521662 522498 557106 522734
rect 557342 522498 557426 522734
rect 557662 522498 589182 522734
rect 589418 522498 589502 522734
rect 589738 522498 592650 522734
rect -8726 522414 592650 522498
rect -8726 522178 -5814 522414
rect -5578 522178 -5494 522414
rect -5258 522178 17106 522414
rect 17342 522178 17426 522414
rect 17662 522178 53106 522414
rect 53342 522178 53426 522414
rect 53662 522178 89106 522414
rect 89342 522178 89426 522414
rect 89662 522178 125106 522414
rect 125342 522178 125426 522414
rect 125662 522178 161106 522414
rect 161342 522178 161426 522414
rect 161662 522178 197106 522414
rect 197342 522178 197426 522414
rect 197662 522178 233106 522414
rect 233342 522178 233426 522414
rect 233662 522178 269106 522414
rect 269342 522178 269426 522414
rect 269662 522178 305106 522414
rect 305342 522178 305426 522414
rect 305662 522178 341106 522414
rect 341342 522178 341426 522414
rect 341662 522178 377106 522414
rect 377342 522178 377426 522414
rect 377662 522178 413106 522414
rect 413342 522178 413426 522414
rect 413662 522178 449106 522414
rect 449342 522178 449426 522414
rect 449662 522178 485106 522414
rect 485342 522178 485426 522414
rect 485662 522178 521106 522414
rect 521342 522178 521426 522414
rect 521662 522178 557106 522414
rect 557342 522178 557426 522414
rect 557662 522178 589182 522414
rect 589418 522178 589502 522414
rect 589738 522178 592650 522414
rect -8726 522146 592650 522178
rect -8726 519014 592650 519046
rect -8726 518778 -4854 519014
rect -4618 518778 -4534 519014
rect -4298 518778 13386 519014
rect 13622 518778 13706 519014
rect 13942 518778 49386 519014
rect 49622 518778 49706 519014
rect 49942 518778 85386 519014
rect 85622 518778 85706 519014
rect 85942 518778 121386 519014
rect 121622 518778 121706 519014
rect 121942 518778 157386 519014
rect 157622 518778 157706 519014
rect 157942 518778 193386 519014
rect 193622 518778 193706 519014
rect 193942 518778 229386 519014
rect 229622 518778 229706 519014
rect 229942 518778 265386 519014
rect 265622 518778 265706 519014
rect 265942 518778 301386 519014
rect 301622 518778 301706 519014
rect 301942 518778 337386 519014
rect 337622 518778 337706 519014
rect 337942 518778 373386 519014
rect 373622 518778 373706 519014
rect 373942 518778 409386 519014
rect 409622 518778 409706 519014
rect 409942 518778 445386 519014
rect 445622 518778 445706 519014
rect 445942 518778 481386 519014
rect 481622 518778 481706 519014
rect 481942 518778 517386 519014
rect 517622 518778 517706 519014
rect 517942 518778 553386 519014
rect 553622 518778 553706 519014
rect 553942 518778 588222 519014
rect 588458 518778 588542 519014
rect 588778 518778 592650 519014
rect -8726 518694 592650 518778
rect -8726 518458 -4854 518694
rect -4618 518458 -4534 518694
rect -4298 518458 13386 518694
rect 13622 518458 13706 518694
rect 13942 518458 49386 518694
rect 49622 518458 49706 518694
rect 49942 518458 85386 518694
rect 85622 518458 85706 518694
rect 85942 518458 121386 518694
rect 121622 518458 121706 518694
rect 121942 518458 157386 518694
rect 157622 518458 157706 518694
rect 157942 518458 193386 518694
rect 193622 518458 193706 518694
rect 193942 518458 229386 518694
rect 229622 518458 229706 518694
rect 229942 518458 265386 518694
rect 265622 518458 265706 518694
rect 265942 518458 301386 518694
rect 301622 518458 301706 518694
rect 301942 518458 337386 518694
rect 337622 518458 337706 518694
rect 337942 518458 373386 518694
rect 373622 518458 373706 518694
rect 373942 518458 409386 518694
rect 409622 518458 409706 518694
rect 409942 518458 445386 518694
rect 445622 518458 445706 518694
rect 445942 518458 481386 518694
rect 481622 518458 481706 518694
rect 481942 518458 517386 518694
rect 517622 518458 517706 518694
rect 517942 518458 553386 518694
rect 553622 518458 553706 518694
rect 553942 518458 588222 518694
rect 588458 518458 588542 518694
rect 588778 518458 592650 518694
rect -8726 518426 592650 518458
rect -8726 515294 592650 515326
rect -8726 515058 -3894 515294
rect -3658 515058 -3574 515294
rect -3338 515058 9666 515294
rect 9902 515058 9986 515294
rect 10222 515058 45666 515294
rect 45902 515058 45986 515294
rect 46222 515058 81666 515294
rect 81902 515058 81986 515294
rect 82222 515058 117666 515294
rect 117902 515058 117986 515294
rect 118222 515058 153666 515294
rect 153902 515058 153986 515294
rect 154222 515058 189666 515294
rect 189902 515058 189986 515294
rect 190222 515058 225666 515294
rect 225902 515058 225986 515294
rect 226222 515058 261666 515294
rect 261902 515058 261986 515294
rect 262222 515058 297666 515294
rect 297902 515058 297986 515294
rect 298222 515058 333666 515294
rect 333902 515058 333986 515294
rect 334222 515058 369666 515294
rect 369902 515058 369986 515294
rect 370222 515058 405666 515294
rect 405902 515058 405986 515294
rect 406222 515058 441666 515294
rect 441902 515058 441986 515294
rect 442222 515058 477666 515294
rect 477902 515058 477986 515294
rect 478222 515058 513666 515294
rect 513902 515058 513986 515294
rect 514222 515058 549666 515294
rect 549902 515058 549986 515294
rect 550222 515058 587262 515294
rect 587498 515058 587582 515294
rect 587818 515058 592650 515294
rect -8726 514974 592650 515058
rect -8726 514738 -3894 514974
rect -3658 514738 -3574 514974
rect -3338 514738 9666 514974
rect 9902 514738 9986 514974
rect 10222 514738 45666 514974
rect 45902 514738 45986 514974
rect 46222 514738 81666 514974
rect 81902 514738 81986 514974
rect 82222 514738 117666 514974
rect 117902 514738 117986 514974
rect 118222 514738 153666 514974
rect 153902 514738 153986 514974
rect 154222 514738 189666 514974
rect 189902 514738 189986 514974
rect 190222 514738 225666 514974
rect 225902 514738 225986 514974
rect 226222 514738 261666 514974
rect 261902 514738 261986 514974
rect 262222 514738 297666 514974
rect 297902 514738 297986 514974
rect 298222 514738 333666 514974
rect 333902 514738 333986 514974
rect 334222 514738 369666 514974
rect 369902 514738 369986 514974
rect 370222 514738 405666 514974
rect 405902 514738 405986 514974
rect 406222 514738 441666 514974
rect 441902 514738 441986 514974
rect 442222 514738 477666 514974
rect 477902 514738 477986 514974
rect 478222 514738 513666 514974
rect 513902 514738 513986 514974
rect 514222 514738 549666 514974
rect 549902 514738 549986 514974
rect 550222 514738 587262 514974
rect 587498 514738 587582 514974
rect 587818 514738 592650 514974
rect -8726 514706 592650 514738
rect -8726 511574 592650 511606
rect -8726 511338 -2934 511574
rect -2698 511338 -2614 511574
rect -2378 511338 5946 511574
rect 6182 511338 6266 511574
rect 6502 511338 41946 511574
rect 42182 511338 42266 511574
rect 42502 511338 77946 511574
rect 78182 511338 78266 511574
rect 78502 511338 113946 511574
rect 114182 511338 114266 511574
rect 114502 511338 149946 511574
rect 150182 511338 150266 511574
rect 150502 511338 185946 511574
rect 186182 511338 186266 511574
rect 186502 511338 221946 511574
rect 222182 511338 222266 511574
rect 222502 511338 257946 511574
rect 258182 511338 258266 511574
rect 258502 511338 293946 511574
rect 294182 511338 294266 511574
rect 294502 511338 329946 511574
rect 330182 511338 330266 511574
rect 330502 511338 365946 511574
rect 366182 511338 366266 511574
rect 366502 511338 401946 511574
rect 402182 511338 402266 511574
rect 402502 511338 437946 511574
rect 438182 511338 438266 511574
rect 438502 511338 473946 511574
rect 474182 511338 474266 511574
rect 474502 511338 509946 511574
rect 510182 511338 510266 511574
rect 510502 511338 545946 511574
rect 546182 511338 546266 511574
rect 546502 511338 581946 511574
rect 582182 511338 582266 511574
rect 582502 511338 586302 511574
rect 586538 511338 586622 511574
rect 586858 511338 592650 511574
rect -8726 511254 592650 511338
rect -8726 511018 -2934 511254
rect -2698 511018 -2614 511254
rect -2378 511018 5946 511254
rect 6182 511018 6266 511254
rect 6502 511018 41946 511254
rect 42182 511018 42266 511254
rect 42502 511018 77946 511254
rect 78182 511018 78266 511254
rect 78502 511018 113946 511254
rect 114182 511018 114266 511254
rect 114502 511018 149946 511254
rect 150182 511018 150266 511254
rect 150502 511018 185946 511254
rect 186182 511018 186266 511254
rect 186502 511018 221946 511254
rect 222182 511018 222266 511254
rect 222502 511018 257946 511254
rect 258182 511018 258266 511254
rect 258502 511018 293946 511254
rect 294182 511018 294266 511254
rect 294502 511018 329946 511254
rect 330182 511018 330266 511254
rect 330502 511018 365946 511254
rect 366182 511018 366266 511254
rect 366502 511018 401946 511254
rect 402182 511018 402266 511254
rect 402502 511018 437946 511254
rect 438182 511018 438266 511254
rect 438502 511018 473946 511254
rect 474182 511018 474266 511254
rect 474502 511018 509946 511254
rect 510182 511018 510266 511254
rect 510502 511018 545946 511254
rect 546182 511018 546266 511254
rect 546502 511018 581946 511254
rect 582182 511018 582266 511254
rect 582502 511018 586302 511254
rect 586538 511018 586622 511254
rect 586858 511018 592650 511254
rect -8726 510986 592650 511018
rect -8726 507854 592650 507886
rect -8726 507618 -1974 507854
rect -1738 507618 -1654 507854
rect -1418 507618 2226 507854
rect 2462 507618 2546 507854
rect 2782 507618 38226 507854
rect 38462 507618 38546 507854
rect 38782 507618 74226 507854
rect 74462 507618 74546 507854
rect 74782 507618 110226 507854
rect 110462 507618 110546 507854
rect 110782 507618 146226 507854
rect 146462 507618 146546 507854
rect 146782 507618 182226 507854
rect 182462 507618 182546 507854
rect 182782 507618 218226 507854
rect 218462 507618 218546 507854
rect 218782 507618 254226 507854
rect 254462 507618 254546 507854
rect 254782 507618 290226 507854
rect 290462 507618 290546 507854
rect 290782 507618 326226 507854
rect 326462 507618 326546 507854
rect 326782 507618 362226 507854
rect 362462 507618 362546 507854
rect 362782 507618 398226 507854
rect 398462 507618 398546 507854
rect 398782 507618 434226 507854
rect 434462 507618 434546 507854
rect 434782 507618 470226 507854
rect 470462 507618 470546 507854
rect 470782 507618 506226 507854
rect 506462 507618 506546 507854
rect 506782 507618 542226 507854
rect 542462 507618 542546 507854
rect 542782 507618 578226 507854
rect 578462 507618 578546 507854
rect 578782 507618 585342 507854
rect 585578 507618 585662 507854
rect 585898 507618 592650 507854
rect -8726 507534 592650 507618
rect -8726 507298 -1974 507534
rect -1738 507298 -1654 507534
rect -1418 507298 2226 507534
rect 2462 507298 2546 507534
rect 2782 507298 38226 507534
rect 38462 507298 38546 507534
rect 38782 507298 74226 507534
rect 74462 507298 74546 507534
rect 74782 507298 110226 507534
rect 110462 507298 110546 507534
rect 110782 507298 146226 507534
rect 146462 507298 146546 507534
rect 146782 507298 182226 507534
rect 182462 507298 182546 507534
rect 182782 507298 218226 507534
rect 218462 507298 218546 507534
rect 218782 507298 254226 507534
rect 254462 507298 254546 507534
rect 254782 507298 290226 507534
rect 290462 507298 290546 507534
rect 290782 507298 326226 507534
rect 326462 507298 326546 507534
rect 326782 507298 362226 507534
rect 362462 507298 362546 507534
rect 362782 507298 398226 507534
rect 398462 507298 398546 507534
rect 398782 507298 434226 507534
rect 434462 507298 434546 507534
rect 434782 507298 470226 507534
rect 470462 507298 470546 507534
rect 470782 507298 506226 507534
rect 506462 507298 506546 507534
rect 506782 507298 542226 507534
rect 542462 507298 542546 507534
rect 542782 507298 578226 507534
rect 578462 507298 578546 507534
rect 578782 507298 585342 507534
rect 585578 507298 585662 507534
rect 585898 507298 592650 507534
rect -8726 507266 592650 507298
rect -8726 497894 592650 497926
rect -8726 497658 -8694 497894
rect -8458 497658 -8374 497894
rect -8138 497658 28266 497894
rect 28502 497658 28586 497894
rect 28822 497658 64266 497894
rect 64502 497658 64586 497894
rect 64822 497658 100266 497894
rect 100502 497658 100586 497894
rect 100822 497658 136266 497894
rect 136502 497658 136586 497894
rect 136822 497658 172266 497894
rect 172502 497658 172586 497894
rect 172822 497658 208266 497894
rect 208502 497658 208586 497894
rect 208822 497658 244266 497894
rect 244502 497658 244586 497894
rect 244822 497658 280266 497894
rect 280502 497658 280586 497894
rect 280822 497658 316266 497894
rect 316502 497658 316586 497894
rect 316822 497658 352266 497894
rect 352502 497658 352586 497894
rect 352822 497658 388266 497894
rect 388502 497658 388586 497894
rect 388822 497658 424266 497894
rect 424502 497658 424586 497894
rect 424822 497658 460266 497894
rect 460502 497658 460586 497894
rect 460822 497658 496266 497894
rect 496502 497658 496586 497894
rect 496822 497658 532266 497894
rect 532502 497658 532586 497894
rect 532822 497658 568266 497894
rect 568502 497658 568586 497894
rect 568822 497658 592062 497894
rect 592298 497658 592382 497894
rect 592618 497658 592650 497894
rect -8726 497574 592650 497658
rect -8726 497338 -8694 497574
rect -8458 497338 -8374 497574
rect -8138 497338 28266 497574
rect 28502 497338 28586 497574
rect 28822 497338 64266 497574
rect 64502 497338 64586 497574
rect 64822 497338 100266 497574
rect 100502 497338 100586 497574
rect 100822 497338 136266 497574
rect 136502 497338 136586 497574
rect 136822 497338 172266 497574
rect 172502 497338 172586 497574
rect 172822 497338 208266 497574
rect 208502 497338 208586 497574
rect 208822 497338 244266 497574
rect 244502 497338 244586 497574
rect 244822 497338 280266 497574
rect 280502 497338 280586 497574
rect 280822 497338 316266 497574
rect 316502 497338 316586 497574
rect 316822 497338 352266 497574
rect 352502 497338 352586 497574
rect 352822 497338 388266 497574
rect 388502 497338 388586 497574
rect 388822 497338 424266 497574
rect 424502 497338 424586 497574
rect 424822 497338 460266 497574
rect 460502 497338 460586 497574
rect 460822 497338 496266 497574
rect 496502 497338 496586 497574
rect 496822 497338 532266 497574
rect 532502 497338 532586 497574
rect 532822 497338 568266 497574
rect 568502 497338 568586 497574
rect 568822 497338 592062 497574
rect 592298 497338 592382 497574
rect 592618 497338 592650 497574
rect -8726 497306 592650 497338
rect -8726 494174 592650 494206
rect -8726 493938 -7734 494174
rect -7498 493938 -7414 494174
rect -7178 493938 24546 494174
rect 24782 493938 24866 494174
rect 25102 493938 60546 494174
rect 60782 493938 60866 494174
rect 61102 493938 96546 494174
rect 96782 493938 96866 494174
rect 97102 493938 132546 494174
rect 132782 493938 132866 494174
rect 133102 493938 168546 494174
rect 168782 493938 168866 494174
rect 169102 493938 204546 494174
rect 204782 493938 204866 494174
rect 205102 493938 240546 494174
rect 240782 493938 240866 494174
rect 241102 493938 276546 494174
rect 276782 493938 276866 494174
rect 277102 493938 312546 494174
rect 312782 493938 312866 494174
rect 313102 493938 348546 494174
rect 348782 493938 348866 494174
rect 349102 493938 384546 494174
rect 384782 493938 384866 494174
rect 385102 493938 420546 494174
rect 420782 493938 420866 494174
rect 421102 493938 456546 494174
rect 456782 493938 456866 494174
rect 457102 493938 492546 494174
rect 492782 493938 492866 494174
rect 493102 493938 528546 494174
rect 528782 493938 528866 494174
rect 529102 493938 564546 494174
rect 564782 493938 564866 494174
rect 565102 493938 591102 494174
rect 591338 493938 591422 494174
rect 591658 493938 592650 494174
rect -8726 493854 592650 493938
rect -8726 493618 -7734 493854
rect -7498 493618 -7414 493854
rect -7178 493618 24546 493854
rect 24782 493618 24866 493854
rect 25102 493618 60546 493854
rect 60782 493618 60866 493854
rect 61102 493618 96546 493854
rect 96782 493618 96866 493854
rect 97102 493618 132546 493854
rect 132782 493618 132866 493854
rect 133102 493618 168546 493854
rect 168782 493618 168866 493854
rect 169102 493618 204546 493854
rect 204782 493618 204866 493854
rect 205102 493618 240546 493854
rect 240782 493618 240866 493854
rect 241102 493618 276546 493854
rect 276782 493618 276866 493854
rect 277102 493618 312546 493854
rect 312782 493618 312866 493854
rect 313102 493618 348546 493854
rect 348782 493618 348866 493854
rect 349102 493618 384546 493854
rect 384782 493618 384866 493854
rect 385102 493618 420546 493854
rect 420782 493618 420866 493854
rect 421102 493618 456546 493854
rect 456782 493618 456866 493854
rect 457102 493618 492546 493854
rect 492782 493618 492866 493854
rect 493102 493618 528546 493854
rect 528782 493618 528866 493854
rect 529102 493618 564546 493854
rect 564782 493618 564866 493854
rect 565102 493618 591102 493854
rect 591338 493618 591422 493854
rect 591658 493618 592650 493854
rect -8726 493586 592650 493618
rect -8726 490454 592650 490486
rect -8726 490218 -6774 490454
rect -6538 490218 -6454 490454
rect -6218 490218 20826 490454
rect 21062 490218 21146 490454
rect 21382 490218 56826 490454
rect 57062 490218 57146 490454
rect 57382 490218 92826 490454
rect 93062 490218 93146 490454
rect 93382 490218 128826 490454
rect 129062 490218 129146 490454
rect 129382 490218 164826 490454
rect 165062 490218 165146 490454
rect 165382 490218 200826 490454
rect 201062 490218 201146 490454
rect 201382 490218 236826 490454
rect 237062 490218 237146 490454
rect 237382 490218 272826 490454
rect 273062 490218 273146 490454
rect 273382 490218 308826 490454
rect 309062 490218 309146 490454
rect 309382 490218 344826 490454
rect 345062 490218 345146 490454
rect 345382 490218 380826 490454
rect 381062 490218 381146 490454
rect 381382 490218 416826 490454
rect 417062 490218 417146 490454
rect 417382 490218 452826 490454
rect 453062 490218 453146 490454
rect 453382 490218 488826 490454
rect 489062 490218 489146 490454
rect 489382 490218 524826 490454
rect 525062 490218 525146 490454
rect 525382 490218 560826 490454
rect 561062 490218 561146 490454
rect 561382 490218 590142 490454
rect 590378 490218 590462 490454
rect 590698 490218 592650 490454
rect -8726 490134 592650 490218
rect -8726 489898 -6774 490134
rect -6538 489898 -6454 490134
rect -6218 489898 20826 490134
rect 21062 489898 21146 490134
rect 21382 489898 56826 490134
rect 57062 489898 57146 490134
rect 57382 489898 92826 490134
rect 93062 489898 93146 490134
rect 93382 489898 128826 490134
rect 129062 489898 129146 490134
rect 129382 489898 164826 490134
rect 165062 489898 165146 490134
rect 165382 489898 200826 490134
rect 201062 489898 201146 490134
rect 201382 489898 236826 490134
rect 237062 489898 237146 490134
rect 237382 489898 272826 490134
rect 273062 489898 273146 490134
rect 273382 489898 308826 490134
rect 309062 489898 309146 490134
rect 309382 489898 344826 490134
rect 345062 489898 345146 490134
rect 345382 489898 380826 490134
rect 381062 489898 381146 490134
rect 381382 489898 416826 490134
rect 417062 489898 417146 490134
rect 417382 489898 452826 490134
rect 453062 489898 453146 490134
rect 453382 489898 488826 490134
rect 489062 489898 489146 490134
rect 489382 489898 524826 490134
rect 525062 489898 525146 490134
rect 525382 489898 560826 490134
rect 561062 489898 561146 490134
rect 561382 489898 590142 490134
rect 590378 489898 590462 490134
rect 590698 489898 592650 490134
rect -8726 489866 592650 489898
rect -8726 486734 592650 486766
rect -8726 486498 -5814 486734
rect -5578 486498 -5494 486734
rect -5258 486498 17106 486734
rect 17342 486498 17426 486734
rect 17662 486498 53106 486734
rect 53342 486498 53426 486734
rect 53662 486498 89106 486734
rect 89342 486498 89426 486734
rect 89662 486498 125106 486734
rect 125342 486498 125426 486734
rect 125662 486498 161106 486734
rect 161342 486498 161426 486734
rect 161662 486498 197106 486734
rect 197342 486498 197426 486734
rect 197662 486498 233106 486734
rect 233342 486498 233426 486734
rect 233662 486498 269106 486734
rect 269342 486498 269426 486734
rect 269662 486498 305106 486734
rect 305342 486498 305426 486734
rect 305662 486498 341106 486734
rect 341342 486498 341426 486734
rect 341662 486498 377106 486734
rect 377342 486498 377426 486734
rect 377662 486498 413106 486734
rect 413342 486498 413426 486734
rect 413662 486498 449106 486734
rect 449342 486498 449426 486734
rect 449662 486498 485106 486734
rect 485342 486498 485426 486734
rect 485662 486498 521106 486734
rect 521342 486498 521426 486734
rect 521662 486498 557106 486734
rect 557342 486498 557426 486734
rect 557662 486498 589182 486734
rect 589418 486498 589502 486734
rect 589738 486498 592650 486734
rect -8726 486414 592650 486498
rect -8726 486178 -5814 486414
rect -5578 486178 -5494 486414
rect -5258 486178 17106 486414
rect 17342 486178 17426 486414
rect 17662 486178 53106 486414
rect 53342 486178 53426 486414
rect 53662 486178 89106 486414
rect 89342 486178 89426 486414
rect 89662 486178 125106 486414
rect 125342 486178 125426 486414
rect 125662 486178 161106 486414
rect 161342 486178 161426 486414
rect 161662 486178 197106 486414
rect 197342 486178 197426 486414
rect 197662 486178 233106 486414
rect 233342 486178 233426 486414
rect 233662 486178 269106 486414
rect 269342 486178 269426 486414
rect 269662 486178 305106 486414
rect 305342 486178 305426 486414
rect 305662 486178 341106 486414
rect 341342 486178 341426 486414
rect 341662 486178 377106 486414
rect 377342 486178 377426 486414
rect 377662 486178 413106 486414
rect 413342 486178 413426 486414
rect 413662 486178 449106 486414
rect 449342 486178 449426 486414
rect 449662 486178 485106 486414
rect 485342 486178 485426 486414
rect 485662 486178 521106 486414
rect 521342 486178 521426 486414
rect 521662 486178 557106 486414
rect 557342 486178 557426 486414
rect 557662 486178 589182 486414
rect 589418 486178 589502 486414
rect 589738 486178 592650 486414
rect -8726 486146 592650 486178
rect -8726 483014 592650 483046
rect -8726 482778 -4854 483014
rect -4618 482778 -4534 483014
rect -4298 482778 13386 483014
rect 13622 482778 13706 483014
rect 13942 482778 49386 483014
rect 49622 482778 49706 483014
rect 49942 482778 85386 483014
rect 85622 482778 85706 483014
rect 85942 482778 121386 483014
rect 121622 482778 121706 483014
rect 121942 482778 157386 483014
rect 157622 482778 157706 483014
rect 157942 482778 193386 483014
rect 193622 482778 193706 483014
rect 193942 482778 229386 483014
rect 229622 482778 229706 483014
rect 229942 482778 265386 483014
rect 265622 482778 265706 483014
rect 265942 482778 301386 483014
rect 301622 482778 301706 483014
rect 301942 482778 337386 483014
rect 337622 482778 337706 483014
rect 337942 482778 373386 483014
rect 373622 482778 373706 483014
rect 373942 482778 409386 483014
rect 409622 482778 409706 483014
rect 409942 482778 445386 483014
rect 445622 482778 445706 483014
rect 445942 482778 481386 483014
rect 481622 482778 481706 483014
rect 481942 482778 517386 483014
rect 517622 482778 517706 483014
rect 517942 482778 553386 483014
rect 553622 482778 553706 483014
rect 553942 482778 588222 483014
rect 588458 482778 588542 483014
rect 588778 482778 592650 483014
rect -8726 482694 592650 482778
rect -8726 482458 -4854 482694
rect -4618 482458 -4534 482694
rect -4298 482458 13386 482694
rect 13622 482458 13706 482694
rect 13942 482458 49386 482694
rect 49622 482458 49706 482694
rect 49942 482458 85386 482694
rect 85622 482458 85706 482694
rect 85942 482458 121386 482694
rect 121622 482458 121706 482694
rect 121942 482458 157386 482694
rect 157622 482458 157706 482694
rect 157942 482458 193386 482694
rect 193622 482458 193706 482694
rect 193942 482458 229386 482694
rect 229622 482458 229706 482694
rect 229942 482458 265386 482694
rect 265622 482458 265706 482694
rect 265942 482458 301386 482694
rect 301622 482458 301706 482694
rect 301942 482458 337386 482694
rect 337622 482458 337706 482694
rect 337942 482458 373386 482694
rect 373622 482458 373706 482694
rect 373942 482458 409386 482694
rect 409622 482458 409706 482694
rect 409942 482458 445386 482694
rect 445622 482458 445706 482694
rect 445942 482458 481386 482694
rect 481622 482458 481706 482694
rect 481942 482458 517386 482694
rect 517622 482458 517706 482694
rect 517942 482458 553386 482694
rect 553622 482458 553706 482694
rect 553942 482458 588222 482694
rect 588458 482458 588542 482694
rect 588778 482458 592650 482694
rect -8726 482426 592650 482458
rect -8726 479294 592650 479326
rect -8726 479058 -3894 479294
rect -3658 479058 -3574 479294
rect -3338 479058 9666 479294
rect 9902 479058 9986 479294
rect 10222 479058 45666 479294
rect 45902 479058 45986 479294
rect 46222 479058 81666 479294
rect 81902 479058 81986 479294
rect 82222 479058 117666 479294
rect 117902 479058 117986 479294
rect 118222 479058 153666 479294
rect 153902 479058 153986 479294
rect 154222 479058 189666 479294
rect 189902 479058 189986 479294
rect 190222 479058 225666 479294
rect 225902 479058 225986 479294
rect 226222 479058 261666 479294
rect 261902 479058 261986 479294
rect 262222 479058 297666 479294
rect 297902 479058 297986 479294
rect 298222 479058 333666 479294
rect 333902 479058 333986 479294
rect 334222 479058 369666 479294
rect 369902 479058 369986 479294
rect 370222 479058 405666 479294
rect 405902 479058 405986 479294
rect 406222 479058 441666 479294
rect 441902 479058 441986 479294
rect 442222 479058 477666 479294
rect 477902 479058 477986 479294
rect 478222 479058 513666 479294
rect 513902 479058 513986 479294
rect 514222 479058 549666 479294
rect 549902 479058 549986 479294
rect 550222 479058 587262 479294
rect 587498 479058 587582 479294
rect 587818 479058 592650 479294
rect -8726 478974 592650 479058
rect -8726 478738 -3894 478974
rect -3658 478738 -3574 478974
rect -3338 478738 9666 478974
rect 9902 478738 9986 478974
rect 10222 478738 45666 478974
rect 45902 478738 45986 478974
rect 46222 478738 81666 478974
rect 81902 478738 81986 478974
rect 82222 478738 117666 478974
rect 117902 478738 117986 478974
rect 118222 478738 153666 478974
rect 153902 478738 153986 478974
rect 154222 478738 189666 478974
rect 189902 478738 189986 478974
rect 190222 478738 225666 478974
rect 225902 478738 225986 478974
rect 226222 478738 261666 478974
rect 261902 478738 261986 478974
rect 262222 478738 297666 478974
rect 297902 478738 297986 478974
rect 298222 478738 333666 478974
rect 333902 478738 333986 478974
rect 334222 478738 369666 478974
rect 369902 478738 369986 478974
rect 370222 478738 405666 478974
rect 405902 478738 405986 478974
rect 406222 478738 441666 478974
rect 441902 478738 441986 478974
rect 442222 478738 477666 478974
rect 477902 478738 477986 478974
rect 478222 478738 513666 478974
rect 513902 478738 513986 478974
rect 514222 478738 549666 478974
rect 549902 478738 549986 478974
rect 550222 478738 587262 478974
rect 587498 478738 587582 478974
rect 587818 478738 592650 478974
rect -8726 478706 592650 478738
rect -8726 475574 592650 475606
rect -8726 475338 -2934 475574
rect -2698 475338 -2614 475574
rect -2378 475338 5946 475574
rect 6182 475338 6266 475574
rect 6502 475338 41946 475574
rect 42182 475338 42266 475574
rect 42502 475338 77946 475574
rect 78182 475338 78266 475574
rect 78502 475338 113946 475574
rect 114182 475338 114266 475574
rect 114502 475338 149946 475574
rect 150182 475338 150266 475574
rect 150502 475338 185946 475574
rect 186182 475338 186266 475574
rect 186502 475338 221946 475574
rect 222182 475338 222266 475574
rect 222502 475338 257946 475574
rect 258182 475338 258266 475574
rect 258502 475338 293946 475574
rect 294182 475338 294266 475574
rect 294502 475338 329946 475574
rect 330182 475338 330266 475574
rect 330502 475338 365946 475574
rect 366182 475338 366266 475574
rect 366502 475338 401946 475574
rect 402182 475338 402266 475574
rect 402502 475338 437946 475574
rect 438182 475338 438266 475574
rect 438502 475338 473946 475574
rect 474182 475338 474266 475574
rect 474502 475338 509946 475574
rect 510182 475338 510266 475574
rect 510502 475338 545946 475574
rect 546182 475338 546266 475574
rect 546502 475338 581946 475574
rect 582182 475338 582266 475574
rect 582502 475338 586302 475574
rect 586538 475338 586622 475574
rect 586858 475338 592650 475574
rect -8726 475254 592650 475338
rect -8726 475018 -2934 475254
rect -2698 475018 -2614 475254
rect -2378 475018 5946 475254
rect 6182 475018 6266 475254
rect 6502 475018 41946 475254
rect 42182 475018 42266 475254
rect 42502 475018 77946 475254
rect 78182 475018 78266 475254
rect 78502 475018 113946 475254
rect 114182 475018 114266 475254
rect 114502 475018 149946 475254
rect 150182 475018 150266 475254
rect 150502 475018 185946 475254
rect 186182 475018 186266 475254
rect 186502 475018 221946 475254
rect 222182 475018 222266 475254
rect 222502 475018 257946 475254
rect 258182 475018 258266 475254
rect 258502 475018 293946 475254
rect 294182 475018 294266 475254
rect 294502 475018 329946 475254
rect 330182 475018 330266 475254
rect 330502 475018 365946 475254
rect 366182 475018 366266 475254
rect 366502 475018 401946 475254
rect 402182 475018 402266 475254
rect 402502 475018 437946 475254
rect 438182 475018 438266 475254
rect 438502 475018 473946 475254
rect 474182 475018 474266 475254
rect 474502 475018 509946 475254
rect 510182 475018 510266 475254
rect 510502 475018 545946 475254
rect 546182 475018 546266 475254
rect 546502 475018 581946 475254
rect 582182 475018 582266 475254
rect 582502 475018 586302 475254
rect 586538 475018 586622 475254
rect 586858 475018 592650 475254
rect -8726 474986 592650 475018
rect -8726 471854 592650 471886
rect -8726 471618 -1974 471854
rect -1738 471618 -1654 471854
rect -1418 471618 2226 471854
rect 2462 471618 2546 471854
rect 2782 471618 38226 471854
rect 38462 471618 38546 471854
rect 38782 471618 74226 471854
rect 74462 471618 74546 471854
rect 74782 471618 110226 471854
rect 110462 471618 110546 471854
rect 110782 471618 146226 471854
rect 146462 471618 146546 471854
rect 146782 471618 182226 471854
rect 182462 471618 182546 471854
rect 182782 471618 218226 471854
rect 218462 471618 218546 471854
rect 218782 471618 254226 471854
rect 254462 471618 254546 471854
rect 254782 471618 290226 471854
rect 290462 471618 290546 471854
rect 290782 471618 326226 471854
rect 326462 471618 326546 471854
rect 326782 471618 362226 471854
rect 362462 471618 362546 471854
rect 362782 471618 398226 471854
rect 398462 471618 398546 471854
rect 398782 471618 434226 471854
rect 434462 471618 434546 471854
rect 434782 471618 470226 471854
rect 470462 471618 470546 471854
rect 470782 471618 506226 471854
rect 506462 471618 506546 471854
rect 506782 471618 542226 471854
rect 542462 471618 542546 471854
rect 542782 471618 578226 471854
rect 578462 471618 578546 471854
rect 578782 471618 585342 471854
rect 585578 471618 585662 471854
rect 585898 471618 592650 471854
rect -8726 471534 592650 471618
rect -8726 471298 -1974 471534
rect -1738 471298 -1654 471534
rect -1418 471298 2226 471534
rect 2462 471298 2546 471534
rect 2782 471298 38226 471534
rect 38462 471298 38546 471534
rect 38782 471298 74226 471534
rect 74462 471298 74546 471534
rect 74782 471298 110226 471534
rect 110462 471298 110546 471534
rect 110782 471298 146226 471534
rect 146462 471298 146546 471534
rect 146782 471298 182226 471534
rect 182462 471298 182546 471534
rect 182782 471298 218226 471534
rect 218462 471298 218546 471534
rect 218782 471298 254226 471534
rect 254462 471298 254546 471534
rect 254782 471298 290226 471534
rect 290462 471298 290546 471534
rect 290782 471298 326226 471534
rect 326462 471298 326546 471534
rect 326782 471298 362226 471534
rect 362462 471298 362546 471534
rect 362782 471298 398226 471534
rect 398462 471298 398546 471534
rect 398782 471298 434226 471534
rect 434462 471298 434546 471534
rect 434782 471298 470226 471534
rect 470462 471298 470546 471534
rect 470782 471298 506226 471534
rect 506462 471298 506546 471534
rect 506782 471298 542226 471534
rect 542462 471298 542546 471534
rect 542782 471298 578226 471534
rect 578462 471298 578546 471534
rect 578782 471298 585342 471534
rect 585578 471298 585662 471534
rect 585898 471298 592650 471534
rect -8726 471266 592650 471298
rect -8726 461894 592650 461926
rect -8726 461658 -8694 461894
rect -8458 461658 -8374 461894
rect -8138 461658 28266 461894
rect 28502 461658 28586 461894
rect 28822 461658 64266 461894
rect 64502 461658 64586 461894
rect 64822 461658 100266 461894
rect 100502 461658 100586 461894
rect 100822 461658 136266 461894
rect 136502 461658 136586 461894
rect 136822 461658 172266 461894
rect 172502 461658 172586 461894
rect 172822 461658 208266 461894
rect 208502 461658 208586 461894
rect 208822 461658 244266 461894
rect 244502 461658 244586 461894
rect 244822 461658 280266 461894
rect 280502 461658 280586 461894
rect 280822 461658 316266 461894
rect 316502 461658 316586 461894
rect 316822 461658 352266 461894
rect 352502 461658 352586 461894
rect 352822 461658 388266 461894
rect 388502 461658 388586 461894
rect 388822 461658 424266 461894
rect 424502 461658 424586 461894
rect 424822 461658 460266 461894
rect 460502 461658 460586 461894
rect 460822 461658 496266 461894
rect 496502 461658 496586 461894
rect 496822 461658 532266 461894
rect 532502 461658 532586 461894
rect 532822 461658 568266 461894
rect 568502 461658 568586 461894
rect 568822 461658 592062 461894
rect 592298 461658 592382 461894
rect 592618 461658 592650 461894
rect -8726 461574 592650 461658
rect -8726 461338 -8694 461574
rect -8458 461338 -8374 461574
rect -8138 461338 28266 461574
rect 28502 461338 28586 461574
rect 28822 461338 64266 461574
rect 64502 461338 64586 461574
rect 64822 461338 100266 461574
rect 100502 461338 100586 461574
rect 100822 461338 136266 461574
rect 136502 461338 136586 461574
rect 136822 461338 172266 461574
rect 172502 461338 172586 461574
rect 172822 461338 208266 461574
rect 208502 461338 208586 461574
rect 208822 461338 244266 461574
rect 244502 461338 244586 461574
rect 244822 461338 280266 461574
rect 280502 461338 280586 461574
rect 280822 461338 316266 461574
rect 316502 461338 316586 461574
rect 316822 461338 352266 461574
rect 352502 461338 352586 461574
rect 352822 461338 388266 461574
rect 388502 461338 388586 461574
rect 388822 461338 424266 461574
rect 424502 461338 424586 461574
rect 424822 461338 460266 461574
rect 460502 461338 460586 461574
rect 460822 461338 496266 461574
rect 496502 461338 496586 461574
rect 496822 461338 532266 461574
rect 532502 461338 532586 461574
rect 532822 461338 568266 461574
rect 568502 461338 568586 461574
rect 568822 461338 592062 461574
rect 592298 461338 592382 461574
rect 592618 461338 592650 461574
rect -8726 461306 592650 461338
rect -8726 458174 592650 458206
rect -8726 457938 -7734 458174
rect -7498 457938 -7414 458174
rect -7178 457938 24546 458174
rect 24782 457938 24866 458174
rect 25102 457938 60546 458174
rect 60782 457938 60866 458174
rect 61102 457938 96546 458174
rect 96782 457938 96866 458174
rect 97102 457938 132546 458174
rect 132782 457938 132866 458174
rect 133102 457938 168546 458174
rect 168782 457938 168866 458174
rect 169102 457938 204546 458174
rect 204782 457938 204866 458174
rect 205102 457938 240546 458174
rect 240782 457938 240866 458174
rect 241102 457938 276546 458174
rect 276782 457938 276866 458174
rect 277102 457938 312546 458174
rect 312782 457938 312866 458174
rect 313102 457938 348546 458174
rect 348782 457938 348866 458174
rect 349102 457938 384546 458174
rect 384782 457938 384866 458174
rect 385102 457938 420546 458174
rect 420782 457938 420866 458174
rect 421102 457938 456546 458174
rect 456782 457938 456866 458174
rect 457102 457938 492546 458174
rect 492782 457938 492866 458174
rect 493102 457938 528546 458174
rect 528782 457938 528866 458174
rect 529102 457938 564546 458174
rect 564782 457938 564866 458174
rect 565102 457938 591102 458174
rect 591338 457938 591422 458174
rect 591658 457938 592650 458174
rect -8726 457854 592650 457938
rect -8726 457618 -7734 457854
rect -7498 457618 -7414 457854
rect -7178 457618 24546 457854
rect 24782 457618 24866 457854
rect 25102 457618 60546 457854
rect 60782 457618 60866 457854
rect 61102 457618 96546 457854
rect 96782 457618 96866 457854
rect 97102 457618 132546 457854
rect 132782 457618 132866 457854
rect 133102 457618 168546 457854
rect 168782 457618 168866 457854
rect 169102 457618 204546 457854
rect 204782 457618 204866 457854
rect 205102 457618 240546 457854
rect 240782 457618 240866 457854
rect 241102 457618 276546 457854
rect 276782 457618 276866 457854
rect 277102 457618 312546 457854
rect 312782 457618 312866 457854
rect 313102 457618 348546 457854
rect 348782 457618 348866 457854
rect 349102 457618 384546 457854
rect 384782 457618 384866 457854
rect 385102 457618 420546 457854
rect 420782 457618 420866 457854
rect 421102 457618 456546 457854
rect 456782 457618 456866 457854
rect 457102 457618 492546 457854
rect 492782 457618 492866 457854
rect 493102 457618 528546 457854
rect 528782 457618 528866 457854
rect 529102 457618 564546 457854
rect 564782 457618 564866 457854
rect 565102 457618 591102 457854
rect 591338 457618 591422 457854
rect 591658 457618 592650 457854
rect -8726 457586 592650 457618
rect -8726 454454 592650 454486
rect -8726 454218 -6774 454454
rect -6538 454218 -6454 454454
rect -6218 454218 20826 454454
rect 21062 454218 21146 454454
rect 21382 454218 56826 454454
rect 57062 454218 57146 454454
rect 57382 454218 92826 454454
rect 93062 454218 93146 454454
rect 93382 454218 128826 454454
rect 129062 454218 129146 454454
rect 129382 454218 164826 454454
rect 165062 454218 165146 454454
rect 165382 454218 200826 454454
rect 201062 454218 201146 454454
rect 201382 454218 236826 454454
rect 237062 454218 237146 454454
rect 237382 454218 272826 454454
rect 273062 454218 273146 454454
rect 273382 454218 308826 454454
rect 309062 454218 309146 454454
rect 309382 454218 344826 454454
rect 345062 454218 345146 454454
rect 345382 454218 380826 454454
rect 381062 454218 381146 454454
rect 381382 454218 416826 454454
rect 417062 454218 417146 454454
rect 417382 454218 452826 454454
rect 453062 454218 453146 454454
rect 453382 454218 488826 454454
rect 489062 454218 489146 454454
rect 489382 454218 524826 454454
rect 525062 454218 525146 454454
rect 525382 454218 560826 454454
rect 561062 454218 561146 454454
rect 561382 454218 590142 454454
rect 590378 454218 590462 454454
rect 590698 454218 592650 454454
rect -8726 454134 592650 454218
rect -8726 453898 -6774 454134
rect -6538 453898 -6454 454134
rect -6218 453898 20826 454134
rect 21062 453898 21146 454134
rect 21382 453898 56826 454134
rect 57062 453898 57146 454134
rect 57382 453898 92826 454134
rect 93062 453898 93146 454134
rect 93382 453898 128826 454134
rect 129062 453898 129146 454134
rect 129382 453898 164826 454134
rect 165062 453898 165146 454134
rect 165382 453898 200826 454134
rect 201062 453898 201146 454134
rect 201382 453898 236826 454134
rect 237062 453898 237146 454134
rect 237382 453898 272826 454134
rect 273062 453898 273146 454134
rect 273382 453898 308826 454134
rect 309062 453898 309146 454134
rect 309382 453898 344826 454134
rect 345062 453898 345146 454134
rect 345382 453898 380826 454134
rect 381062 453898 381146 454134
rect 381382 453898 416826 454134
rect 417062 453898 417146 454134
rect 417382 453898 452826 454134
rect 453062 453898 453146 454134
rect 453382 453898 488826 454134
rect 489062 453898 489146 454134
rect 489382 453898 524826 454134
rect 525062 453898 525146 454134
rect 525382 453898 560826 454134
rect 561062 453898 561146 454134
rect 561382 453898 590142 454134
rect 590378 453898 590462 454134
rect 590698 453898 592650 454134
rect -8726 453866 592650 453898
rect -8726 450734 592650 450766
rect -8726 450498 -5814 450734
rect -5578 450498 -5494 450734
rect -5258 450498 17106 450734
rect 17342 450498 17426 450734
rect 17662 450498 53106 450734
rect 53342 450498 53426 450734
rect 53662 450498 89106 450734
rect 89342 450498 89426 450734
rect 89662 450498 125106 450734
rect 125342 450498 125426 450734
rect 125662 450498 161106 450734
rect 161342 450498 161426 450734
rect 161662 450498 197106 450734
rect 197342 450498 197426 450734
rect 197662 450498 233106 450734
rect 233342 450498 233426 450734
rect 233662 450498 269106 450734
rect 269342 450498 269426 450734
rect 269662 450498 305106 450734
rect 305342 450498 305426 450734
rect 305662 450498 341106 450734
rect 341342 450498 341426 450734
rect 341662 450498 377106 450734
rect 377342 450498 377426 450734
rect 377662 450498 413106 450734
rect 413342 450498 413426 450734
rect 413662 450498 449106 450734
rect 449342 450498 449426 450734
rect 449662 450498 485106 450734
rect 485342 450498 485426 450734
rect 485662 450498 521106 450734
rect 521342 450498 521426 450734
rect 521662 450498 557106 450734
rect 557342 450498 557426 450734
rect 557662 450498 589182 450734
rect 589418 450498 589502 450734
rect 589738 450498 592650 450734
rect -8726 450414 592650 450498
rect -8726 450178 -5814 450414
rect -5578 450178 -5494 450414
rect -5258 450178 17106 450414
rect 17342 450178 17426 450414
rect 17662 450178 53106 450414
rect 53342 450178 53426 450414
rect 53662 450178 89106 450414
rect 89342 450178 89426 450414
rect 89662 450178 125106 450414
rect 125342 450178 125426 450414
rect 125662 450178 161106 450414
rect 161342 450178 161426 450414
rect 161662 450178 197106 450414
rect 197342 450178 197426 450414
rect 197662 450178 233106 450414
rect 233342 450178 233426 450414
rect 233662 450178 269106 450414
rect 269342 450178 269426 450414
rect 269662 450178 305106 450414
rect 305342 450178 305426 450414
rect 305662 450178 341106 450414
rect 341342 450178 341426 450414
rect 341662 450178 377106 450414
rect 377342 450178 377426 450414
rect 377662 450178 413106 450414
rect 413342 450178 413426 450414
rect 413662 450178 449106 450414
rect 449342 450178 449426 450414
rect 449662 450178 485106 450414
rect 485342 450178 485426 450414
rect 485662 450178 521106 450414
rect 521342 450178 521426 450414
rect 521662 450178 557106 450414
rect 557342 450178 557426 450414
rect 557662 450178 589182 450414
rect 589418 450178 589502 450414
rect 589738 450178 592650 450414
rect -8726 450146 592650 450178
rect -8726 447014 592650 447046
rect -8726 446778 -4854 447014
rect -4618 446778 -4534 447014
rect -4298 446778 13386 447014
rect 13622 446778 13706 447014
rect 13942 446778 49386 447014
rect 49622 446778 49706 447014
rect 49942 446778 85386 447014
rect 85622 446778 85706 447014
rect 85942 446778 121386 447014
rect 121622 446778 121706 447014
rect 121942 446778 157386 447014
rect 157622 446778 157706 447014
rect 157942 446778 193386 447014
rect 193622 446778 193706 447014
rect 193942 446778 229386 447014
rect 229622 446778 229706 447014
rect 229942 446778 265386 447014
rect 265622 446778 265706 447014
rect 265942 446778 301386 447014
rect 301622 446778 301706 447014
rect 301942 446778 337386 447014
rect 337622 446778 337706 447014
rect 337942 446778 373386 447014
rect 373622 446778 373706 447014
rect 373942 446778 409386 447014
rect 409622 446778 409706 447014
rect 409942 446778 445386 447014
rect 445622 446778 445706 447014
rect 445942 446778 481386 447014
rect 481622 446778 481706 447014
rect 481942 446778 517386 447014
rect 517622 446778 517706 447014
rect 517942 446778 553386 447014
rect 553622 446778 553706 447014
rect 553942 446778 588222 447014
rect 588458 446778 588542 447014
rect 588778 446778 592650 447014
rect -8726 446694 592650 446778
rect -8726 446458 -4854 446694
rect -4618 446458 -4534 446694
rect -4298 446458 13386 446694
rect 13622 446458 13706 446694
rect 13942 446458 49386 446694
rect 49622 446458 49706 446694
rect 49942 446458 85386 446694
rect 85622 446458 85706 446694
rect 85942 446458 121386 446694
rect 121622 446458 121706 446694
rect 121942 446458 157386 446694
rect 157622 446458 157706 446694
rect 157942 446458 193386 446694
rect 193622 446458 193706 446694
rect 193942 446458 229386 446694
rect 229622 446458 229706 446694
rect 229942 446458 265386 446694
rect 265622 446458 265706 446694
rect 265942 446458 301386 446694
rect 301622 446458 301706 446694
rect 301942 446458 337386 446694
rect 337622 446458 337706 446694
rect 337942 446458 373386 446694
rect 373622 446458 373706 446694
rect 373942 446458 409386 446694
rect 409622 446458 409706 446694
rect 409942 446458 445386 446694
rect 445622 446458 445706 446694
rect 445942 446458 481386 446694
rect 481622 446458 481706 446694
rect 481942 446458 517386 446694
rect 517622 446458 517706 446694
rect 517942 446458 553386 446694
rect 553622 446458 553706 446694
rect 553942 446458 588222 446694
rect 588458 446458 588542 446694
rect 588778 446458 592650 446694
rect -8726 446426 592650 446458
rect -8726 443294 592650 443326
rect -8726 443058 -3894 443294
rect -3658 443058 -3574 443294
rect -3338 443058 9666 443294
rect 9902 443058 9986 443294
rect 10222 443058 45666 443294
rect 45902 443058 45986 443294
rect 46222 443058 81666 443294
rect 81902 443058 81986 443294
rect 82222 443058 117666 443294
rect 117902 443058 117986 443294
rect 118222 443058 153666 443294
rect 153902 443058 153986 443294
rect 154222 443058 189666 443294
rect 189902 443058 189986 443294
rect 190222 443058 225666 443294
rect 225902 443058 225986 443294
rect 226222 443058 261666 443294
rect 261902 443058 261986 443294
rect 262222 443058 297666 443294
rect 297902 443058 297986 443294
rect 298222 443058 333666 443294
rect 333902 443058 333986 443294
rect 334222 443058 369666 443294
rect 369902 443058 369986 443294
rect 370222 443058 405666 443294
rect 405902 443058 405986 443294
rect 406222 443058 441666 443294
rect 441902 443058 441986 443294
rect 442222 443058 477666 443294
rect 477902 443058 477986 443294
rect 478222 443058 513666 443294
rect 513902 443058 513986 443294
rect 514222 443058 549666 443294
rect 549902 443058 549986 443294
rect 550222 443058 587262 443294
rect 587498 443058 587582 443294
rect 587818 443058 592650 443294
rect -8726 442974 592650 443058
rect -8726 442738 -3894 442974
rect -3658 442738 -3574 442974
rect -3338 442738 9666 442974
rect 9902 442738 9986 442974
rect 10222 442738 45666 442974
rect 45902 442738 45986 442974
rect 46222 442738 81666 442974
rect 81902 442738 81986 442974
rect 82222 442738 117666 442974
rect 117902 442738 117986 442974
rect 118222 442738 153666 442974
rect 153902 442738 153986 442974
rect 154222 442738 189666 442974
rect 189902 442738 189986 442974
rect 190222 442738 225666 442974
rect 225902 442738 225986 442974
rect 226222 442738 261666 442974
rect 261902 442738 261986 442974
rect 262222 442738 297666 442974
rect 297902 442738 297986 442974
rect 298222 442738 333666 442974
rect 333902 442738 333986 442974
rect 334222 442738 369666 442974
rect 369902 442738 369986 442974
rect 370222 442738 405666 442974
rect 405902 442738 405986 442974
rect 406222 442738 441666 442974
rect 441902 442738 441986 442974
rect 442222 442738 477666 442974
rect 477902 442738 477986 442974
rect 478222 442738 513666 442974
rect 513902 442738 513986 442974
rect 514222 442738 549666 442974
rect 549902 442738 549986 442974
rect 550222 442738 587262 442974
rect 587498 442738 587582 442974
rect 587818 442738 592650 442974
rect -8726 442706 592650 442738
rect -8726 439574 592650 439606
rect -8726 439338 -2934 439574
rect -2698 439338 -2614 439574
rect -2378 439338 5946 439574
rect 6182 439338 6266 439574
rect 6502 439338 41946 439574
rect 42182 439338 42266 439574
rect 42502 439338 77946 439574
rect 78182 439338 78266 439574
rect 78502 439338 113946 439574
rect 114182 439338 114266 439574
rect 114502 439338 149946 439574
rect 150182 439338 150266 439574
rect 150502 439338 185946 439574
rect 186182 439338 186266 439574
rect 186502 439338 221946 439574
rect 222182 439338 222266 439574
rect 222502 439338 257946 439574
rect 258182 439338 258266 439574
rect 258502 439338 293946 439574
rect 294182 439338 294266 439574
rect 294502 439338 329946 439574
rect 330182 439338 330266 439574
rect 330502 439338 365946 439574
rect 366182 439338 366266 439574
rect 366502 439338 401946 439574
rect 402182 439338 402266 439574
rect 402502 439338 437946 439574
rect 438182 439338 438266 439574
rect 438502 439338 473946 439574
rect 474182 439338 474266 439574
rect 474502 439338 509946 439574
rect 510182 439338 510266 439574
rect 510502 439338 545946 439574
rect 546182 439338 546266 439574
rect 546502 439338 581946 439574
rect 582182 439338 582266 439574
rect 582502 439338 586302 439574
rect 586538 439338 586622 439574
rect 586858 439338 592650 439574
rect -8726 439254 592650 439338
rect -8726 439018 -2934 439254
rect -2698 439018 -2614 439254
rect -2378 439018 5946 439254
rect 6182 439018 6266 439254
rect 6502 439018 41946 439254
rect 42182 439018 42266 439254
rect 42502 439018 77946 439254
rect 78182 439018 78266 439254
rect 78502 439018 113946 439254
rect 114182 439018 114266 439254
rect 114502 439018 149946 439254
rect 150182 439018 150266 439254
rect 150502 439018 185946 439254
rect 186182 439018 186266 439254
rect 186502 439018 221946 439254
rect 222182 439018 222266 439254
rect 222502 439018 257946 439254
rect 258182 439018 258266 439254
rect 258502 439018 293946 439254
rect 294182 439018 294266 439254
rect 294502 439018 329946 439254
rect 330182 439018 330266 439254
rect 330502 439018 365946 439254
rect 366182 439018 366266 439254
rect 366502 439018 401946 439254
rect 402182 439018 402266 439254
rect 402502 439018 437946 439254
rect 438182 439018 438266 439254
rect 438502 439018 473946 439254
rect 474182 439018 474266 439254
rect 474502 439018 509946 439254
rect 510182 439018 510266 439254
rect 510502 439018 545946 439254
rect 546182 439018 546266 439254
rect 546502 439018 581946 439254
rect 582182 439018 582266 439254
rect 582502 439018 586302 439254
rect 586538 439018 586622 439254
rect 586858 439018 592650 439254
rect -8726 438986 592650 439018
rect -8726 435854 592650 435886
rect -8726 435618 -1974 435854
rect -1738 435618 -1654 435854
rect -1418 435618 2226 435854
rect 2462 435618 2546 435854
rect 2782 435618 38226 435854
rect 38462 435618 38546 435854
rect 38782 435618 74226 435854
rect 74462 435618 74546 435854
rect 74782 435618 110226 435854
rect 110462 435618 110546 435854
rect 110782 435618 146226 435854
rect 146462 435618 146546 435854
rect 146782 435618 182226 435854
rect 182462 435618 182546 435854
rect 182782 435618 218226 435854
rect 218462 435618 218546 435854
rect 218782 435618 254226 435854
rect 254462 435618 254546 435854
rect 254782 435618 290226 435854
rect 290462 435618 290546 435854
rect 290782 435618 326226 435854
rect 326462 435618 326546 435854
rect 326782 435618 362226 435854
rect 362462 435618 362546 435854
rect 362782 435618 398226 435854
rect 398462 435618 398546 435854
rect 398782 435618 434226 435854
rect 434462 435618 434546 435854
rect 434782 435618 470226 435854
rect 470462 435618 470546 435854
rect 470782 435618 506226 435854
rect 506462 435618 506546 435854
rect 506782 435618 542226 435854
rect 542462 435618 542546 435854
rect 542782 435618 578226 435854
rect 578462 435618 578546 435854
rect 578782 435618 585342 435854
rect 585578 435618 585662 435854
rect 585898 435618 592650 435854
rect -8726 435534 592650 435618
rect -8726 435298 -1974 435534
rect -1738 435298 -1654 435534
rect -1418 435298 2226 435534
rect 2462 435298 2546 435534
rect 2782 435298 38226 435534
rect 38462 435298 38546 435534
rect 38782 435298 74226 435534
rect 74462 435298 74546 435534
rect 74782 435298 110226 435534
rect 110462 435298 110546 435534
rect 110782 435298 146226 435534
rect 146462 435298 146546 435534
rect 146782 435298 182226 435534
rect 182462 435298 182546 435534
rect 182782 435298 218226 435534
rect 218462 435298 218546 435534
rect 218782 435298 254226 435534
rect 254462 435298 254546 435534
rect 254782 435298 290226 435534
rect 290462 435298 290546 435534
rect 290782 435298 326226 435534
rect 326462 435298 326546 435534
rect 326782 435298 362226 435534
rect 362462 435298 362546 435534
rect 362782 435298 398226 435534
rect 398462 435298 398546 435534
rect 398782 435298 434226 435534
rect 434462 435298 434546 435534
rect 434782 435298 470226 435534
rect 470462 435298 470546 435534
rect 470782 435298 506226 435534
rect 506462 435298 506546 435534
rect 506782 435298 542226 435534
rect 542462 435298 542546 435534
rect 542782 435298 578226 435534
rect 578462 435298 578546 435534
rect 578782 435298 585342 435534
rect 585578 435298 585662 435534
rect 585898 435298 592650 435534
rect -8726 435266 592650 435298
rect -8726 425894 592650 425926
rect -8726 425658 -8694 425894
rect -8458 425658 -8374 425894
rect -8138 425658 28266 425894
rect 28502 425658 28586 425894
rect 28822 425658 64266 425894
rect 64502 425658 64586 425894
rect 64822 425658 100266 425894
rect 100502 425658 100586 425894
rect 100822 425658 136266 425894
rect 136502 425658 136586 425894
rect 136822 425658 172266 425894
rect 172502 425658 172586 425894
rect 172822 425658 208266 425894
rect 208502 425658 208586 425894
rect 208822 425658 244266 425894
rect 244502 425658 244586 425894
rect 244822 425658 280266 425894
rect 280502 425658 280586 425894
rect 280822 425658 316266 425894
rect 316502 425658 316586 425894
rect 316822 425658 352266 425894
rect 352502 425658 352586 425894
rect 352822 425658 388266 425894
rect 388502 425658 388586 425894
rect 388822 425658 424266 425894
rect 424502 425658 424586 425894
rect 424822 425658 460266 425894
rect 460502 425658 460586 425894
rect 460822 425658 496266 425894
rect 496502 425658 496586 425894
rect 496822 425658 532266 425894
rect 532502 425658 532586 425894
rect 532822 425658 568266 425894
rect 568502 425658 568586 425894
rect 568822 425658 592062 425894
rect 592298 425658 592382 425894
rect 592618 425658 592650 425894
rect -8726 425574 592650 425658
rect -8726 425338 -8694 425574
rect -8458 425338 -8374 425574
rect -8138 425338 28266 425574
rect 28502 425338 28586 425574
rect 28822 425338 64266 425574
rect 64502 425338 64586 425574
rect 64822 425338 100266 425574
rect 100502 425338 100586 425574
rect 100822 425338 136266 425574
rect 136502 425338 136586 425574
rect 136822 425338 172266 425574
rect 172502 425338 172586 425574
rect 172822 425338 208266 425574
rect 208502 425338 208586 425574
rect 208822 425338 244266 425574
rect 244502 425338 244586 425574
rect 244822 425338 280266 425574
rect 280502 425338 280586 425574
rect 280822 425338 316266 425574
rect 316502 425338 316586 425574
rect 316822 425338 352266 425574
rect 352502 425338 352586 425574
rect 352822 425338 388266 425574
rect 388502 425338 388586 425574
rect 388822 425338 424266 425574
rect 424502 425338 424586 425574
rect 424822 425338 460266 425574
rect 460502 425338 460586 425574
rect 460822 425338 496266 425574
rect 496502 425338 496586 425574
rect 496822 425338 532266 425574
rect 532502 425338 532586 425574
rect 532822 425338 568266 425574
rect 568502 425338 568586 425574
rect 568822 425338 592062 425574
rect 592298 425338 592382 425574
rect 592618 425338 592650 425574
rect -8726 425306 592650 425338
rect -8726 422174 592650 422206
rect -8726 421938 -7734 422174
rect -7498 421938 -7414 422174
rect -7178 421938 24546 422174
rect 24782 421938 24866 422174
rect 25102 421938 60546 422174
rect 60782 421938 60866 422174
rect 61102 421938 96546 422174
rect 96782 421938 96866 422174
rect 97102 421938 132546 422174
rect 132782 421938 132866 422174
rect 133102 421938 168546 422174
rect 168782 421938 168866 422174
rect 169102 421938 204546 422174
rect 204782 421938 204866 422174
rect 205102 421938 240546 422174
rect 240782 421938 240866 422174
rect 241102 421938 276546 422174
rect 276782 421938 276866 422174
rect 277102 421938 312546 422174
rect 312782 421938 312866 422174
rect 313102 421938 348546 422174
rect 348782 421938 348866 422174
rect 349102 421938 384546 422174
rect 384782 421938 384866 422174
rect 385102 421938 420546 422174
rect 420782 421938 420866 422174
rect 421102 421938 456546 422174
rect 456782 421938 456866 422174
rect 457102 421938 492546 422174
rect 492782 421938 492866 422174
rect 493102 421938 528546 422174
rect 528782 421938 528866 422174
rect 529102 421938 564546 422174
rect 564782 421938 564866 422174
rect 565102 421938 591102 422174
rect 591338 421938 591422 422174
rect 591658 421938 592650 422174
rect -8726 421854 592650 421938
rect -8726 421618 -7734 421854
rect -7498 421618 -7414 421854
rect -7178 421618 24546 421854
rect 24782 421618 24866 421854
rect 25102 421618 60546 421854
rect 60782 421618 60866 421854
rect 61102 421618 96546 421854
rect 96782 421618 96866 421854
rect 97102 421618 132546 421854
rect 132782 421618 132866 421854
rect 133102 421618 168546 421854
rect 168782 421618 168866 421854
rect 169102 421618 204546 421854
rect 204782 421618 204866 421854
rect 205102 421618 240546 421854
rect 240782 421618 240866 421854
rect 241102 421618 276546 421854
rect 276782 421618 276866 421854
rect 277102 421618 312546 421854
rect 312782 421618 312866 421854
rect 313102 421618 348546 421854
rect 348782 421618 348866 421854
rect 349102 421618 384546 421854
rect 384782 421618 384866 421854
rect 385102 421618 420546 421854
rect 420782 421618 420866 421854
rect 421102 421618 456546 421854
rect 456782 421618 456866 421854
rect 457102 421618 492546 421854
rect 492782 421618 492866 421854
rect 493102 421618 528546 421854
rect 528782 421618 528866 421854
rect 529102 421618 564546 421854
rect 564782 421618 564866 421854
rect 565102 421618 591102 421854
rect 591338 421618 591422 421854
rect 591658 421618 592650 421854
rect -8726 421586 592650 421618
rect -8726 418454 592650 418486
rect -8726 418218 -6774 418454
rect -6538 418218 -6454 418454
rect -6218 418218 20826 418454
rect 21062 418218 21146 418454
rect 21382 418218 56826 418454
rect 57062 418218 57146 418454
rect 57382 418218 92826 418454
rect 93062 418218 93146 418454
rect 93382 418218 128826 418454
rect 129062 418218 129146 418454
rect 129382 418218 164826 418454
rect 165062 418218 165146 418454
rect 165382 418218 200826 418454
rect 201062 418218 201146 418454
rect 201382 418218 236826 418454
rect 237062 418218 237146 418454
rect 237382 418218 272826 418454
rect 273062 418218 273146 418454
rect 273382 418218 308826 418454
rect 309062 418218 309146 418454
rect 309382 418218 344826 418454
rect 345062 418218 345146 418454
rect 345382 418218 380826 418454
rect 381062 418218 381146 418454
rect 381382 418218 416826 418454
rect 417062 418218 417146 418454
rect 417382 418218 452826 418454
rect 453062 418218 453146 418454
rect 453382 418218 488826 418454
rect 489062 418218 489146 418454
rect 489382 418218 524826 418454
rect 525062 418218 525146 418454
rect 525382 418218 560826 418454
rect 561062 418218 561146 418454
rect 561382 418218 590142 418454
rect 590378 418218 590462 418454
rect 590698 418218 592650 418454
rect -8726 418134 592650 418218
rect -8726 417898 -6774 418134
rect -6538 417898 -6454 418134
rect -6218 417898 20826 418134
rect 21062 417898 21146 418134
rect 21382 417898 56826 418134
rect 57062 417898 57146 418134
rect 57382 417898 92826 418134
rect 93062 417898 93146 418134
rect 93382 417898 128826 418134
rect 129062 417898 129146 418134
rect 129382 417898 164826 418134
rect 165062 417898 165146 418134
rect 165382 417898 200826 418134
rect 201062 417898 201146 418134
rect 201382 417898 236826 418134
rect 237062 417898 237146 418134
rect 237382 417898 272826 418134
rect 273062 417898 273146 418134
rect 273382 417898 308826 418134
rect 309062 417898 309146 418134
rect 309382 417898 344826 418134
rect 345062 417898 345146 418134
rect 345382 417898 380826 418134
rect 381062 417898 381146 418134
rect 381382 417898 416826 418134
rect 417062 417898 417146 418134
rect 417382 417898 452826 418134
rect 453062 417898 453146 418134
rect 453382 417898 488826 418134
rect 489062 417898 489146 418134
rect 489382 417898 524826 418134
rect 525062 417898 525146 418134
rect 525382 417898 560826 418134
rect 561062 417898 561146 418134
rect 561382 417898 590142 418134
rect 590378 417898 590462 418134
rect 590698 417898 592650 418134
rect -8726 417866 592650 417898
rect -8726 414734 592650 414766
rect -8726 414498 -5814 414734
rect -5578 414498 -5494 414734
rect -5258 414498 17106 414734
rect 17342 414498 17426 414734
rect 17662 414498 53106 414734
rect 53342 414498 53426 414734
rect 53662 414498 89106 414734
rect 89342 414498 89426 414734
rect 89662 414498 125106 414734
rect 125342 414498 125426 414734
rect 125662 414498 161106 414734
rect 161342 414498 161426 414734
rect 161662 414498 197106 414734
rect 197342 414498 197426 414734
rect 197662 414498 233106 414734
rect 233342 414498 233426 414734
rect 233662 414498 269106 414734
rect 269342 414498 269426 414734
rect 269662 414498 305106 414734
rect 305342 414498 305426 414734
rect 305662 414498 341106 414734
rect 341342 414498 341426 414734
rect 341662 414498 377106 414734
rect 377342 414498 377426 414734
rect 377662 414498 413106 414734
rect 413342 414498 413426 414734
rect 413662 414498 449106 414734
rect 449342 414498 449426 414734
rect 449662 414498 485106 414734
rect 485342 414498 485426 414734
rect 485662 414498 521106 414734
rect 521342 414498 521426 414734
rect 521662 414498 557106 414734
rect 557342 414498 557426 414734
rect 557662 414498 589182 414734
rect 589418 414498 589502 414734
rect 589738 414498 592650 414734
rect -8726 414414 592650 414498
rect -8726 414178 -5814 414414
rect -5578 414178 -5494 414414
rect -5258 414178 17106 414414
rect 17342 414178 17426 414414
rect 17662 414178 53106 414414
rect 53342 414178 53426 414414
rect 53662 414178 89106 414414
rect 89342 414178 89426 414414
rect 89662 414178 125106 414414
rect 125342 414178 125426 414414
rect 125662 414178 161106 414414
rect 161342 414178 161426 414414
rect 161662 414178 197106 414414
rect 197342 414178 197426 414414
rect 197662 414178 233106 414414
rect 233342 414178 233426 414414
rect 233662 414178 269106 414414
rect 269342 414178 269426 414414
rect 269662 414178 305106 414414
rect 305342 414178 305426 414414
rect 305662 414178 341106 414414
rect 341342 414178 341426 414414
rect 341662 414178 377106 414414
rect 377342 414178 377426 414414
rect 377662 414178 413106 414414
rect 413342 414178 413426 414414
rect 413662 414178 449106 414414
rect 449342 414178 449426 414414
rect 449662 414178 485106 414414
rect 485342 414178 485426 414414
rect 485662 414178 521106 414414
rect 521342 414178 521426 414414
rect 521662 414178 557106 414414
rect 557342 414178 557426 414414
rect 557662 414178 589182 414414
rect 589418 414178 589502 414414
rect 589738 414178 592650 414414
rect -8726 414146 592650 414178
rect -8726 411014 592650 411046
rect -8726 410778 -4854 411014
rect -4618 410778 -4534 411014
rect -4298 410778 13386 411014
rect 13622 410778 13706 411014
rect 13942 410778 49386 411014
rect 49622 410778 49706 411014
rect 49942 410778 85386 411014
rect 85622 410778 85706 411014
rect 85942 410778 121386 411014
rect 121622 410778 121706 411014
rect 121942 410778 157386 411014
rect 157622 410778 157706 411014
rect 157942 410778 193386 411014
rect 193622 410778 193706 411014
rect 193942 410778 229386 411014
rect 229622 410778 229706 411014
rect 229942 410778 265386 411014
rect 265622 410778 265706 411014
rect 265942 410778 301386 411014
rect 301622 410778 301706 411014
rect 301942 410778 337386 411014
rect 337622 410778 337706 411014
rect 337942 410778 373386 411014
rect 373622 410778 373706 411014
rect 373942 410778 409386 411014
rect 409622 410778 409706 411014
rect 409942 410778 445386 411014
rect 445622 410778 445706 411014
rect 445942 410778 481386 411014
rect 481622 410778 481706 411014
rect 481942 410778 517386 411014
rect 517622 410778 517706 411014
rect 517942 410778 553386 411014
rect 553622 410778 553706 411014
rect 553942 410778 588222 411014
rect 588458 410778 588542 411014
rect 588778 410778 592650 411014
rect -8726 410694 592650 410778
rect -8726 410458 -4854 410694
rect -4618 410458 -4534 410694
rect -4298 410458 13386 410694
rect 13622 410458 13706 410694
rect 13942 410458 49386 410694
rect 49622 410458 49706 410694
rect 49942 410458 85386 410694
rect 85622 410458 85706 410694
rect 85942 410458 121386 410694
rect 121622 410458 121706 410694
rect 121942 410458 157386 410694
rect 157622 410458 157706 410694
rect 157942 410458 193386 410694
rect 193622 410458 193706 410694
rect 193942 410458 229386 410694
rect 229622 410458 229706 410694
rect 229942 410458 265386 410694
rect 265622 410458 265706 410694
rect 265942 410458 301386 410694
rect 301622 410458 301706 410694
rect 301942 410458 337386 410694
rect 337622 410458 337706 410694
rect 337942 410458 373386 410694
rect 373622 410458 373706 410694
rect 373942 410458 409386 410694
rect 409622 410458 409706 410694
rect 409942 410458 445386 410694
rect 445622 410458 445706 410694
rect 445942 410458 481386 410694
rect 481622 410458 481706 410694
rect 481942 410458 517386 410694
rect 517622 410458 517706 410694
rect 517942 410458 553386 410694
rect 553622 410458 553706 410694
rect 553942 410458 588222 410694
rect 588458 410458 588542 410694
rect 588778 410458 592650 410694
rect -8726 410426 592650 410458
rect -8726 407294 592650 407326
rect -8726 407058 -3894 407294
rect -3658 407058 -3574 407294
rect -3338 407058 9666 407294
rect 9902 407058 9986 407294
rect 10222 407058 45666 407294
rect 45902 407058 45986 407294
rect 46222 407058 81666 407294
rect 81902 407058 81986 407294
rect 82222 407058 117666 407294
rect 117902 407058 117986 407294
rect 118222 407058 153666 407294
rect 153902 407058 153986 407294
rect 154222 407058 189666 407294
rect 189902 407058 189986 407294
rect 190222 407058 225666 407294
rect 225902 407058 225986 407294
rect 226222 407058 261666 407294
rect 261902 407058 261986 407294
rect 262222 407058 297666 407294
rect 297902 407058 297986 407294
rect 298222 407058 333666 407294
rect 333902 407058 333986 407294
rect 334222 407058 369666 407294
rect 369902 407058 369986 407294
rect 370222 407058 405666 407294
rect 405902 407058 405986 407294
rect 406222 407058 441666 407294
rect 441902 407058 441986 407294
rect 442222 407058 477666 407294
rect 477902 407058 477986 407294
rect 478222 407058 513666 407294
rect 513902 407058 513986 407294
rect 514222 407058 549666 407294
rect 549902 407058 549986 407294
rect 550222 407058 587262 407294
rect 587498 407058 587582 407294
rect 587818 407058 592650 407294
rect -8726 406974 592650 407058
rect -8726 406738 -3894 406974
rect -3658 406738 -3574 406974
rect -3338 406738 9666 406974
rect 9902 406738 9986 406974
rect 10222 406738 45666 406974
rect 45902 406738 45986 406974
rect 46222 406738 81666 406974
rect 81902 406738 81986 406974
rect 82222 406738 117666 406974
rect 117902 406738 117986 406974
rect 118222 406738 153666 406974
rect 153902 406738 153986 406974
rect 154222 406738 189666 406974
rect 189902 406738 189986 406974
rect 190222 406738 225666 406974
rect 225902 406738 225986 406974
rect 226222 406738 261666 406974
rect 261902 406738 261986 406974
rect 262222 406738 297666 406974
rect 297902 406738 297986 406974
rect 298222 406738 333666 406974
rect 333902 406738 333986 406974
rect 334222 406738 369666 406974
rect 369902 406738 369986 406974
rect 370222 406738 405666 406974
rect 405902 406738 405986 406974
rect 406222 406738 441666 406974
rect 441902 406738 441986 406974
rect 442222 406738 477666 406974
rect 477902 406738 477986 406974
rect 478222 406738 513666 406974
rect 513902 406738 513986 406974
rect 514222 406738 549666 406974
rect 549902 406738 549986 406974
rect 550222 406738 587262 406974
rect 587498 406738 587582 406974
rect 587818 406738 592650 406974
rect -8726 406706 592650 406738
rect -8726 403574 592650 403606
rect -8726 403338 -2934 403574
rect -2698 403338 -2614 403574
rect -2378 403338 5946 403574
rect 6182 403338 6266 403574
rect 6502 403338 41946 403574
rect 42182 403338 42266 403574
rect 42502 403338 77946 403574
rect 78182 403338 78266 403574
rect 78502 403338 113946 403574
rect 114182 403338 114266 403574
rect 114502 403338 149946 403574
rect 150182 403338 150266 403574
rect 150502 403338 185946 403574
rect 186182 403338 186266 403574
rect 186502 403338 221946 403574
rect 222182 403338 222266 403574
rect 222502 403338 257946 403574
rect 258182 403338 258266 403574
rect 258502 403338 293946 403574
rect 294182 403338 294266 403574
rect 294502 403338 329946 403574
rect 330182 403338 330266 403574
rect 330502 403338 365946 403574
rect 366182 403338 366266 403574
rect 366502 403338 401946 403574
rect 402182 403338 402266 403574
rect 402502 403338 437946 403574
rect 438182 403338 438266 403574
rect 438502 403338 473946 403574
rect 474182 403338 474266 403574
rect 474502 403338 509946 403574
rect 510182 403338 510266 403574
rect 510502 403338 545946 403574
rect 546182 403338 546266 403574
rect 546502 403338 581946 403574
rect 582182 403338 582266 403574
rect 582502 403338 586302 403574
rect 586538 403338 586622 403574
rect 586858 403338 592650 403574
rect -8726 403254 592650 403338
rect -8726 403018 -2934 403254
rect -2698 403018 -2614 403254
rect -2378 403018 5946 403254
rect 6182 403018 6266 403254
rect 6502 403018 41946 403254
rect 42182 403018 42266 403254
rect 42502 403018 77946 403254
rect 78182 403018 78266 403254
rect 78502 403018 113946 403254
rect 114182 403018 114266 403254
rect 114502 403018 149946 403254
rect 150182 403018 150266 403254
rect 150502 403018 185946 403254
rect 186182 403018 186266 403254
rect 186502 403018 221946 403254
rect 222182 403018 222266 403254
rect 222502 403018 257946 403254
rect 258182 403018 258266 403254
rect 258502 403018 293946 403254
rect 294182 403018 294266 403254
rect 294502 403018 329946 403254
rect 330182 403018 330266 403254
rect 330502 403018 365946 403254
rect 366182 403018 366266 403254
rect 366502 403018 401946 403254
rect 402182 403018 402266 403254
rect 402502 403018 437946 403254
rect 438182 403018 438266 403254
rect 438502 403018 473946 403254
rect 474182 403018 474266 403254
rect 474502 403018 509946 403254
rect 510182 403018 510266 403254
rect 510502 403018 545946 403254
rect 546182 403018 546266 403254
rect 546502 403018 581946 403254
rect 582182 403018 582266 403254
rect 582502 403018 586302 403254
rect 586538 403018 586622 403254
rect 586858 403018 592650 403254
rect -8726 402986 592650 403018
rect -8726 399854 592650 399886
rect -8726 399618 -1974 399854
rect -1738 399618 -1654 399854
rect -1418 399618 2226 399854
rect 2462 399618 2546 399854
rect 2782 399618 38226 399854
rect 38462 399618 38546 399854
rect 38782 399618 74226 399854
rect 74462 399618 74546 399854
rect 74782 399618 110226 399854
rect 110462 399618 110546 399854
rect 110782 399618 146226 399854
rect 146462 399618 146546 399854
rect 146782 399618 182226 399854
rect 182462 399618 182546 399854
rect 182782 399618 218226 399854
rect 218462 399618 218546 399854
rect 218782 399618 254226 399854
rect 254462 399618 254546 399854
rect 254782 399618 290226 399854
rect 290462 399618 290546 399854
rect 290782 399618 326226 399854
rect 326462 399618 326546 399854
rect 326782 399618 362226 399854
rect 362462 399618 362546 399854
rect 362782 399618 398226 399854
rect 398462 399618 398546 399854
rect 398782 399618 434226 399854
rect 434462 399618 434546 399854
rect 434782 399618 470226 399854
rect 470462 399618 470546 399854
rect 470782 399618 506226 399854
rect 506462 399618 506546 399854
rect 506782 399618 542226 399854
rect 542462 399618 542546 399854
rect 542782 399618 578226 399854
rect 578462 399618 578546 399854
rect 578782 399618 585342 399854
rect 585578 399618 585662 399854
rect 585898 399618 592650 399854
rect -8726 399534 592650 399618
rect -8726 399298 -1974 399534
rect -1738 399298 -1654 399534
rect -1418 399298 2226 399534
rect 2462 399298 2546 399534
rect 2782 399298 38226 399534
rect 38462 399298 38546 399534
rect 38782 399298 74226 399534
rect 74462 399298 74546 399534
rect 74782 399298 110226 399534
rect 110462 399298 110546 399534
rect 110782 399298 146226 399534
rect 146462 399298 146546 399534
rect 146782 399298 182226 399534
rect 182462 399298 182546 399534
rect 182782 399298 218226 399534
rect 218462 399298 218546 399534
rect 218782 399298 254226 399534
rect 254462 399298 254546 399534
rect 254782 399298 290226 399534
rect 290462 399298 290546 399534
rect 290782 399298 326226 399534
rect 326462 399298 326546 399534
rect 326782 399298 362226 399534
rect 362462 399298 362546 399534
rect 362782 399298 398226 399534
rect 398462 399298 398546 399534
rect 398782 399298 434226 399534
rect 434462 399298 434546 399534
rect 434782 399298 470226 399534
rect 470462 399298 470546 399534
rect 470782 399298 506226 399534
rect 506462 399298 506546 399534
rect 506782 399298 542226 399534
rect 542462 399298 542546 399534
rect 542782 399298 578226 399534
rect 578462 399298 578546 399534
rect 578782 399298 585342 399534
rect 585578 399298 585662 399534
rect 585898 399298 592650 399534
rect -8726 399266 592650 399298
rect -8726 389894 592650 389926
rect -8726 389658 -8694 389894
rect -8458 389658 -8374 389894
rect -8138 389658 28266 389894
rect 28502 389658 28586 389894
rect 28822 389658 64266 389894
rect 64502 389658 64586 389894
rect 64822 389658 100266 389894
rect 100502 389658 100586 389894
rect 100822 389658 136266 389894
rect 136502 389658 136586 389894
rect 136822 389658 172266 389894
rect 172502 389658 172586 389894
rect 172822 389658 208266 389894
rect 208502 389658 208586 389894
rect 208822 389658 244266 389894
rect 244502 389658 244586 389894
rect 244822 389658 280266 389894
rect 280502 389658 280586 389894
rect 280822 389658 316266 389894
rect 316502 389658 316586 389894
rect 316822 389658 352266 389894
rect 352502 389658 352586 389894
rect 352822 389658 388266 389894
rect 388502 389658 388586 389894
rect 388822 389658 424266 389894
rect 424502 389658 424586 389894
rect 424822 389658 460266 389894
rect 460502 389658 460586 389894
rect 460822 389658 496266 389894
rect 496502 389658 496586 389894
rect 496822 389658 532266 389894
rect 532502 389658 532586 389894
rect 532822 389658 568266 389894
rect 568502 389658 568586 389894
rect 568822 389658 592062 389894
rect 592298 389658 592382 389894
rect 592618 389658 592650 389894
rect -8726 389574 592650 389658
rect -8726 389338 -8694 389574
rect -8458 389338 -8374 389574
rect -8138 389338 28266 389574
rect 28502 389338 28586 389574
rect 28822 389338 64266 389574
rect 64502 389338 64586 389574
rect 64822 389338 100266 389574
rect 100502 389338 100586 389574
rect 100822 389338 136266 389574
rect 136502 389338 136586 389574
rect 136822 389338 172266 389574
rect 172502 389338 172586 389574
rect 172822 389338 208266 389574
rect 208502 389338 208586 389574
rect 208822 389338 244266 389574
rect 244502 389338 244586 389574
rect 244822 389338 280266 389574
rect 280502 389338 280586 389574
rect 280822 389338 316266 389574
rect 316502 389338 316586 389574
rect 316822 389338 352266 389574
rect 352502 389338 352586 389574
rect 352822 389338 388266 389574
rect 388502 389338 388586 389574
rect 388822 389338 424266 389574
rect 424502 389338 424586 389574
rect 424822 389338 460266 389574
rect 460502 389338 460586 389574
rect 460822 389338 496266 389574
rect 496502 389338 496586 389574
rect 496822 389338 532266 389574
rect 532502 389338 532586 389574
rect 532822 389338 568266 389574
rect 568502 389338 568586 389574
rect 568822 389338 592062 389574
rect 592298 389338 592382 389574
rect 592618 389338 592650 389574
rect -8726 389306 592650 389338
rect -8726 386174 592650 386206
rect -8726 385938 -7734 386174
rect -7498 385938 -7414 386174
rect -7178 385938 24546 386174
rect 24782 385938 24866 386174
rect 25102 385938 60546 386174
rect 60782 385938 60866 386174
rect 61102 385938 96546 386174
rect 96782 385938 96866 386174
rect 97102 385938 132546 386174
rect 132782 385938 132866 386174
rect 133102 385938 168546 386174
rect 168782 385938 168866 386174
rect 169102 385938 204546 386174
rect 204782 385938 204866 386174
rect 205102 385938 240546 386174
rect 240782 385938 240866 386174
rect 241102 385938 276546 386174
rect 276782 385938 276866 386174
rect 277102 385938 312546 386174
rect 312782 385938 312866 386174
rect 313102 385938 348546 386174
rect 348782 385938 348866 386174
rect 349102 385938 384546 386174
rect 384782 385938 384866 386174
rect 385102 385938 420546 386174
rect 420782 385938 420866 386174
rect 421102 385938 456546 386174
rect 456782 385938 456866 386174
rect 457102 385938 492546 386174
rect 492782 385938 492866 386174
rect 493102 385938 528546 386174
rect 528782 385938 528866 386174
rect 529102 385938 564546 386174
rect 564782 385938 564866 386174
rect 565102 385938 591102 386174
rect 591338 385938 591422 386174
rect 591658 385938 592650 386174
rect -8726 385854 592650 385938
rect -8726 385618 -7734 385854
rect -7498 385618 -7414 385854
rect -7178 385618 24546 385854
rect 24782 385618 24866 385854
rect 25102 385618 60546 385854
rect 60782 385618 60866 385854
rect 61102 385618 96546 385854
rect 96782 385618 96866 385854
rect 97102 385618 132546 385854
rect 132782 385618 132866 385854
rect 133102 385618 168546 385854
rect 168782 385618 168866 385854
rect 169102 385618 204546 385854
rect 204782 385618 204866 385854
rect 205102 385618 240546 385854
rect 240782 385618 240866 385854
rect 241102 385618 276546 385854
rect 276782 385618 276866 385854
rect 277102 385618 312546 385854
rect 312782 385618 312866 385854
rect 313102 385618 348546 385854
rect 348782 385618 348866 385854
rect 349102 385618 384546 385854
rect 384782 385618 384866 385854
rect 385102 385618 420546 385854
rect 420782 385618 420866 385854
rect 421102 385618 456546 385854
rect 456782 385618 456866 385854
rect 457102 385618 492546 385854
rect 492782 385618 492866 385854
rect 493102 385618 528546 385854
rect 528782 385618 528866 385854
rect 529102 385618 564546 385854
rect 564782 385618 564866 385854
rect 565102 385618 591102 385854
rect 591338 385618 591422 385854
rect 591658 385618 592650 385854
rect -8726 385586 592650 385618
rect -8726 382454 592650 382486
rect -8726 382218 -6774 382454
rect -6538 382218 -6454 382454
rect -6218 382218 20826 382454
rect 21062 382218 21146 382454
rect 21382 382218 56826 382454
rect 57062 382218 57146 382454
rect 57382 382218 92826 382454
rect 93062 382218 93146 382454
rect 93382 382218 128826 382454
rect 129062 382218 129146 382454
rect 129382 382218 164826 382454
rect 165062 382218 165146 382454
rect 165382 382218 200826 382454
rect 201062 382218 201146 382454
rect 201382 382218 236826 382454
rect 237062 382218 237146 382454
rect 237382 382218 272826 382454
rect 273062 382218 273146 382454
rect 273382 382218 308826 382454
rect 309062 382218 309146 382454
rect 309382 382218 344826 382454
rect 345062 382218 345146 382454
rect 345382 382218 380826 382454
rect 381062 382218 381146 382454
rect 381382 382218 416826 382454
rect 417062 382218 417146 382454
rect 417382 382218 452826 382454
rect 453062 382218 453146 382454
rect 453382 382218 488826 382454
rect 489062 382218 489146 382454
rect 489382 382218 524826 382454
rect 525062 382218 525146 382454
rect 525382 382218 560826 382454
rect 561062 382218 561146 382454
rect 561382 382218 590142 382454
rect 590378 382218 590462 382454
rect 590698 382218 592650 382454
rect -8726 382134 592650 382218
rect -8726 381898 -6774 382134
rect -6538 381898 -6454 382134
rect -6218 381898 20826 382134
rect 21062 381898 21146 382134
rect 21382 381898 56826 382134
rect 57062 381898 57146 382134
rect 57382 381898 92826 382134
rect 93062 381898 93146 382134
rect 93382 381898 128826 382134
rect 129062 381898 129146 382134
rect 129382 381898 164826 382134
rect 165062 381898 165146 382134
rect 165382 381898 200826 382134
rect 201062 381898 201146 382134
rect 201382 381898 236826 382134
rect 237062 381898 237146 382134
rect 237382 381898 272826 382134
rect 273062 381898 273146 382134
rect 273382 381898 308826 382134
rect 309062 381898 309146 382134
rect 309382 381898 344826 382134
rect 345062 381898 345146 382134
rect 345382 381898 380826 382134
rect 381062 381898 381146 382134
rect 381382 381898 416826 382134
rect 417062 381898 417146 382134
rect 417382 381898 452826 382134
rect 453062 381898 453146 382134
rect 453382 381898 488826 382134
rect 489062 381898 489146 382134
rect 489382 381898 524826 382134
rect 525062 381898 525146 382134
rect 525382 381898 560826 382134
rect 561062 381898 561146 382134
rect 561382 381898 590142 382134
rect 590378 381898 590462 382134
rect 590698 381898 592650 382134
rect -8726 381866 592650 381898
rect -8726 378734 592650 378766
rect -8726 378498 -5814 378734
rect -5578 378498 -5494 378734
rect -5258 378498 17106 378734
rect 17342 378498 17426 378734
rect 17662 378498 53106 378734
rect 53342 378498 53426 378734
rect 53662 378498 89106 378734
rect 89342 378498 89426 378734
rect 89662 378498 125106 378734
rect 125342 378498 125426 378734
rect 125662 378498 161106 378734
rect 161342 378498 161426 378734
rect 161662 378498 197106 378734
rect 197342 378498 197426 378734
rect 197662 378498 233106 378734
rect 233342 378498 233426 378734
rect 233662 378498 269106 378734
rect 269342 378498 269426 378734
rect 269662 378498 305106 378734
rect 305342 378498 305426 378734
rect 305662 378498 341106 378734
rect 341342 378498 341426 378734
rect 341662 378498 377106 378734
rect 377342 378498 377426 378734
rect 377662 378498 413106 378734
rect 413342 378498 413426 378734
rect 413662 378498 449106 378734
rect 449342 378498 449426 378734
rect 449662 378498 485106 378734
rect 485342 378498 485426 378734
rect 485662 378498 521106 378734
rect 521342 378498 521426 378734
rect 521662 378498 557106 378734
rect 557342 378498 557426 378734
rect 557662 378498 589182 378734
rect 589418 378498 589502 378734
rect 589738 378498 592650 378734
rect -8726 378414 592650 378498
rect -8726 378178 -5814 378414
rect -5578 378178 -5494 378414
rect -5258 378178 17106 378414
rect 17342 378178 17426 378414
rect 17662 378178 53106 378414
rect 53342 378178 53426 378414
rect 53662 378178 89106 378414
rect 89342 378178 89426 378414
rect 89662 378178 125106 378414
rect 125342 378178 125426 378414
rect 125662 378178 161106 378414
rect 161342 378178 161426 378414
rect 161662 378178 197106 378414
rect 197342 378178 197426 378414
rect 197662 378178 233106 378414
rect 233342 378178 233426 378414
rect 233662 378178 269106 378414
rect 269342 378178 269426 378414
rect 269662 378178 305106 378414
rect 305342 378178 305426 378414
rect 305662 378178 341106 378414
rect 341342 378178 341426 378414
rect 341662 378178 377106 378414
rect 377342 378178 377426 378414
rect 377662 378178 413106 378414
rect 413342 378178 413426 378414
rect 413662 378178 449106 378414
rect 449342 378178 449426 378414
rect 449662 378178 485106 378414
rect 485342 378178 485426 378414
rect 485662 378178 521106 378414
rect 521342 378178 521426 378414
rect 521662 378178 557106 378414
rect 557342 378178 557426 378414
rect 557662 378178 589182 378414
rect 589418 378178 589502 378414
rect 589738 378178 592650 378414
rect -8726 378146 592650 378178
rect -8726 375014 592650 375046
rect -8726 374778 -4854 375014
rect -4618 374778 -4534 375014
rect -4298 374778 13386 375014
rect 13622 374778 13706 375014
rect 13942 374778 49386 375014
rect 49622 374778 49706 375014
rect 49942 374778 85386 375014
rect 85622 374778 85706 375014
rect 85942 374778 121386 375014
rect 121622 374778 121706 375014
rect 121942 374778 157386 375014
rect 157622 374778 157706 375014
rect 157942 374778 193386 375014
rect 193622 374778 193706 375014
rect 193942 374778 229386 375014
rect 229622 374778 229706 375014
rect 229942 374778 265386 375014
rect 265622 374778 265706 375014
rect 265942 374778 301386 375014
rect 301622 374778 301706 375014
rect 301942 374778 337386 375014
rect 337622 374778 337706 375014
rect 337942 374778 373386 375014
rect 373622 374778 373706 375014
rect 373942 374778 409386 375014
rect 409622 374778 409706 375014
rect 409942 374778 445386 375014
rect 445622 374778 445706 375014
rect 445942 374778 481386 375014
rect 481622 374778 481706 375014
rect 481942 374778 517386 375014
rect 517622 374778 517706 375014
rect 517942 374778 553386 375014
rect 553622 374778 553706 375014
rect 553942 374778 588222 375014
rect 588458 374778 588542 375014
rect 588778 374778 592650 375014
rect -8726 374694 592650 374778
rect -8726 374458 -4854 374694
rect -4618 374458 -4534 374694
rect -4298 374458 13386 374694
rect 13622 374458 13706 374694
rect 13942 374458 49386 374694
rect 49622 374458 49706 374694
rect 49942 374458 85386 374694
rect 85622 374458 85706 374694
rect 85942 374458 121386 374694
rect 121622 374458 121706 374694
rect 121942 374458 157386 374694
rect 157622 374458 157706 374694
rect 157942 374458 193386 374694
rect 193622 374458 193706 374694
rect 193942 374458 229386 374694
rect 229622 374458 229706 374694
rect 229942 374458 265386 374694
rect 265622 374458 265706 374694
rect 265942 374458 301386 374694
rect 301622 374458 301706 374694
rect 301942 374458 337386 374694
rect 337622 374458 337706 374694
rect 337942 374458 373386 374694
rect 373622 374458 373706 374694
rect 373942 374458 409386 374694
rect 409622 374458 409706 374694
rect 409942 374458 445386 374694
rect 445622 374458 445706 374694
rect 445942 374458 481386 374694
rect 481622 374458 481706 374694
rect 481942 374458 517386 374694
rect 517622 374458 517706 374694
rect 517942 374458 553386 374694
rect 553622 374458 553706 374694
rect 553942 374458 588222 374694
rect 588458 374458 588542 374694
rect 588778 374458 592650 374694
rect -8726 374426 592650 374458
rect -8726 371294 592650 371326
rect -8726 371058 -3894 371294
rect -3658 371058 -3574 371294
rect -3338 371058 9666 371294
rect 9902 371058 9986 371294
rect 10222 371058 45666 371294
rect 45902 371058 45986 371294
rect 46222 371058 81666 371294
rect 81902 371058 81986 371294
rect 82222 371058 117666 371294
rect 117902 371058 117986 371294
rect 118222 371058 153666 371294
rect 153902 371058 153986 371294
rect 154222 371058 189666 371294
rect 189902 371058 189986 371294
rect 190222 371058 225666 371294
rect 225902 371058 225986 371294
rect 226222 371058 261666 371294
rect 261902 371058 261986 371294
rect 262222 371058 297666 371294
rect 297902 371058 297986 371294
rect 298222 371058 333666 371294
rect 333902 371058 333986 371294
rect 334222 371058 369666 371294
rect 369902 371058 369986 371294
rect 370222 371058 405666 371294
rect 405902 371058 405986 371294
rect 406222 371058 441666 371294
rect 441902 371058 441986 371294
rect 442222 371058 477666 371294
rect 477902 371058 477986 371294
rect 478222 371058 513666 371294
rect 513902 371058 513986 371294
rect 514222 371058 549666 371294
rect 549902 371058 549986 371294
rect 550222 371058 587262 371294
rect 587498 371058 587582 371294
rect 587818 371058 592650 371294
rect -8726 370974 592650 371058
rect -8726 370738 -3894 370974
rect -3658 370738 -3574 370974
rect -3338 370738 9666 370974
rect 9902 370738 9986 370974
rect 10222 370738 45666 370974
rect 45902 370738 45986 370974
rect 46222 370738 81666 370974
rect 81902 370738 81986 370974
rect 82222 370738 117666 370974
rect 117902 370738 117986 370974
rect 118222 370738 153666 370974
rect 153902 370738 153986 370974
rect 154222 370738 189666 370974
rect 189902 370738 189986 370974
rect 190222 370738 225666 370974
rect 225902 370738 225986 370974
rect 226222 370738 261666 370974
rect 261902 370738 261986 370974
rect 262222 370738 297666 370974
rect 297902 370738 297986 370974
rect 298222 370738 333666 370974
rect 333902 370738 333986 370974
rect 334222 370738 369666 370974
rect 369902 370738 369986 370974
rect 370222 370738 405666 370974
rect 405902 370738 405986 370974
rect 406222 370738 441666 370974
rect 441902 370738 441986 370974
rect 442222 370738 477666 370974
rect 477902 370738 477986 370974
rect 478222 370738 513666 370974
rect 513902 370738 513986 370974
rect 514222 370738 549666 370974
rect 549902 370738 549986 370974
rect 550222 370738 587262 370974
rect 587498 370738 587582 370974
rect 587818 370738 592650 370974
rect -8726 370706 592650 370738
rect -8726 367574 592650 367606
rect -8726 367338 -2934 367574
rect -2698 367338 -2614 367574
rect -2378 367338 5946 367574
rect 6182 367338 6266 367574
rect 6502 367338 41946 367574
rect 42182 367338 42266 367574
rect 42502 367338 77946 367574
rect 78182 367338 78266 367574
rect 78502 367338 113946 367574
rect 114182 367338 114266 367574
rect 114502 367338 149946 367574
rect 150182 367338 150266 367574
rect 150502 367338 185946 367574
rect 186182 367338 186266 367574
rect 186502 367338 221946 367574
rect 222182 367338 222266 367574
rect 222502 367338 257946 367574
rect 258182 367338 258266 367574
rect 258502 367338 293946 367574
rect 294182 367338 294266 367574
rect 294502 367338 329946 367574
rect 330182 367338 330266 367574
rect 330502 367338 365946 367574
rect 366182 367338 366266 367574
rect 366502 367338 401946 367574
rect 402182 367338 402266 367574
rect 402502 367338 437946 367574
rect 438182 367338 438266 367574
rect 438502 367338 473946 367574
rect 474182 367338 474266 367574
rect 474502 367338 509946 367574
rect 510182 367338 510266 367574
rect 510502 367338 545946 367574
rect 546182 367338 546266 367574
rect 546502 367338 581946 367574
rect 582182 367338 582266 367574
rect 582502 367338 586302 367574
rect 586538 367338 586622 367574
rect 586858 367338 592650 367574
rect -8726 367254 592650 367338
rect -8726 367018 -2934 367254
rect -2698 367018 -2614 367254
rect -2378 367018 5946 367254
rect 6182 367018 6266 367254
rect 6502 367018 41946 367254
rect 42182 367018 42266 367254
rect 42502 367018 77946 367254
rect 78182 367018 78266 367254
rect 78502 367018 113946 367254
rect 114182 367018 114266 367254
rect 114502 367018 149946 367254
rect 150182 367018 150266 367254
rect 150502 367018 185946 367254
rect 186182 367018 186266 367254
rect 186502 367018 221946 367254
rect 222182 367018 222266 367254
rect 222502 367018 257946 367254
rect 258182 367018 258266 367254
rect 258502 367018 293946 367254
rect 294182 367018 294266 367254
rect 294502 367018 329946 367254
rect 330182 367018 330266 367254
rect 330502 367018 365946 367254
rect 366182 367018 366266 367254
rect 366502 367018 401946 367254
rect 402182 367018 402266 367254
rect 402502 367018 437946 367254
rect 438182 367018 438266 367254
rect 438502 367018 473946 367254
rect 474182 367018 474266 367254
rect 474502 367018 509946 367254
rect 510182 367018 510266 367254
rect 510502 367018 545946 367254
rect 546182 367018 546266 367254
rect 546502 367018 581946 367254
rect 582182 367018 582266 367254
rect 582502 367018 586302 367254
rect 586538 367018 586622 367254
rect 586858 367018 592650 367254
rect -8726 366986 592650 367018
rect -8726 363854 592650 363886
rect -8726 363618 -1974 363854
rect -1738 363618 -1654 363854
rect -1418 363618 2226 363854
rect 2462 363618 2546 363854
rect 2782 363618 38226 363854
rect 38462 363618 38546 363854
rect 38782 363618 74226 363854
rect 74462 363618 74546 363854
rect 74782 363618 110226 363854
rect 110462 363618 110546 363854
rect 110782 363618 146226 363854
rect 146462 363618 146546 363854
rect 146782 363618 182226 363854
rect 182462 363618 182546 363854
rect 182782 363618 218226 363854
rect 218462 363618 218546 363854
rect 218782 363618 254226 363854
rect 254462 363618 254546 363854
rect 254782 363618 290226 363854
rect 290462 363618 290546 363854
rect 290782 363618 326226 363854
rect 326462 363618 326546 363854
rect 326782 363618 362226 363854
rect 362462 363618 362546 363854
rect 362782 363618 398226 363854
rect 398462 363618 398546 363854
rect 398782 363618 434226 363854
rect 434462 363618 434546 363854
rect 434782 363618 470226 363854
rect 470462 363618 470546 363854
rect 470782 363618 506226 363854
rect 506462 363618 506546 363854
rect 506782 363618 542226 363854
rect 542462 363618 542546 363854
rect 542782 363618 578226 363854
rect 578462 363618 578546 363854
rect 578782 363618 585342 363854
rect 585578 363618 585662 363854
rect 585898 363618 592650 363854
rect -8726 363534 592650 363618
rect -8726 363298 -1974 363534
rect -1738 363298 -1654 363534
rect -1418 363298 2226 363534
rect 2462 363298 2546 363534
rect 2782 363298 38226 363534
rect 38462 363298 38546 363534
rect 38782 363298 74226 363534
rect 74462 363298 74546 363534
rect 74782 363298 110226 363534
rect 110462 363298 110546 363534
rect 110782 363298 146226 363534
rect 146462 363298 146546 363534
rect 146782 363298 182226 363534
rect 182462 363298 182546 363534
rect 182782 363298 218226 363534
rect 218462 363298 218546 363534
rect 218782 363298 254226 363534
rect 254462 363298 254546 363534
rect 254782 363298 290226 363534
rect 290462 363298 290546 363534
rect 290782 363298 326226 363534
rect 326462 363298 326546 363534
rect 326782 363298 362226 363534
rect 362462 363298 362546 363534
rect 362782 363298 398226 363534
rect 398462 363298 398546 363534
rect 398782 363298 434226 363534
rect 434462 363298 434546 363534
rect 434782 363298 470226 363534
rect 470462 363298 470546 363534
rect 470782 363298 506226 363534
rect 506462 363298 506546 363534
rect 506782 363298 542226 363534
rect 542462 363298 542546 363534
rect 542782 363298 578226 363534
rect 578462 363298 578546 363534
rect 578782 363298 585342 363534
rect 585578 363298 585662 363534
rect 585898 363298 592650 363534
rect -8726 363266 592650 363298
rect -8726 353894 592650 353926
rect -8726 353658 -8694 353894
rect -8458 353658 -8374 353894
rect -8138 353658 28266 353894
rect 28502 353658 28586 353894
rect 28822 353658 64266 353894
rect 64502 353658 64586 353894
rect 64822 353658 100266 353894
rect 100502 353658 100586 353894
rect 100822 353658 136266 353894
rect 136502 353658 136586 353894
rect 136822 353658 172266 353894
rect 172502 353658 172586 353894
rect 172822 353658 208266 353894
rect 208502 353658 208586 353894
rect 208822 353658 244266 353894
rect 244502 353658 244586 353894
rect 244822 353658 280266 353894
rect 280502 353658 280586 353894
rect 280822 353658 316266 353894
rect 316502 353658 316586 353894
rect 316822 353658 352266 353894
rect 352502 353658 352586 353894
rect 352822 353658 388266 353894
rect 388502 353658 388586 353894
rect 388822 353658 424266 353894
rect 424502 353658 424586 353894
rect 424822 353658 460266 353894
rect 460502 353658 460586 353894
rect 460822 353658 496266 353894
rect 496502 353658 496586 353894
rect 496822 353658 532266 353894
rect 532502 353658 532586 353894
rect 532822 353658 568266 353894
rect 568502 353658 568586 353894
rect 568822 353658 592062 353894
rect 592298 353658 592382 353894
rect 592618 353658 592650 353894
rect -8726 353574 592650 353658
rect -8726 353338 -8694 353574
rect -8458 353338 -8374 353574
rect -8138 353338 28266 353574
rect 28502 353338 28586 353574
rect 28822 353338 64266 353574
rect 64502 353338 64586 353574
rect 64822 353338 100266 353574
rect 100502 353338 100586 353574
rect 100822 353338 136266 353574
rect 136502 353338 136586 353574
rect 136822 353338 172266 353574
rect 172502 353338 172586 353574
rect 172822 353338 208266 353574
rect 208502 353338 208586 353574
rect 208822 353338 244266 353574
rect 244502 353338 244586 353574
rect 244822 353338 280266 353574
rect 280502 353338 280586 353574
rect 280822 353338 316266 353574
rect 316502 353338 316586 353574
rect 316822 353338 352266 353574
rect 352502 353338 352586 353574
rect 352822 353338 388266 353574
rect 388502 353338 388586 353574
rect 388822 353338 424266 353574
rect 424502 353338 424586 353574
rect 424822 353338 460266 353574
rect 460502 353338 460586 353574
rect 460822 353338 496266 353574
rect 496502 353338 496586 353574
rect 496822 353338 532266 353574
rect 532502 353338 532586 353574
rect 532822 353338 568266 353574
rect 568502 353338 568586 353574
rect 568822 353338 592062 353574
rect 592298 353338 592382 353574
rect 592618 353338 592650 353574
rect -8726 353306 592650 353338
rect -8726 350174 592650 350206
rect -8726 349938 -7734 350174
rect -7498 349938 -7414 350174
rect -7178 349938 24546 350174
rect 24782 349938 24866 350174
rect 25102 349938 60546 350174
rect 60782 349938 60866 350174
rect 61102 349938 96546 350174
rect 96782 349938 96866 350174
rect 97102 349938 132546 350174
rect 132782 349938 132866 350174
rect 133102 349938 168546 350174
rect 168782 349938 168866 350174
rect 169102 349938 204546 350174
rect 204782 349938 204866 350174
rect 205102 349938 240546 350174
rect 240782 349938 240866 350174
rect 241102 349938 276546 350174
rect 276782 349938 276866 350174
rect 277102 349938 312546 350174
rect 312782 349938 312866 350174
rect 313102 349938 348546 350174
rect 348782 349938 348866 350174
rect 349102 349938 384546 350174
rect 384782 349938 384866 350174
rect 385102 349938 420546 350174
rect 420782 349938 420866 350174
rect 421102 349938 456546 350174
rect 456782 349938 456866 350174
rect 457102 349938 492546 350174
rect 492782 349938 492866 350174
rect 493102 349938 528546 350174
rect 528782 349938 528866 350174
rect 529102 349938 564546 350174
rect 564782 349938 564866 350174
rect 565102 349938 591102 350174
rect 591338 349938 591422 350174
rect 591658 349938 592650 350174
rect -8726 349854 592650 349938
rect -8726 349618 -7734 349854
rect -7498 349618 -7414 349854
rect -7178 349618 24546 349854
rect 24782 349618 24866 349854
rect 25102 349618 60546 349854
rect 60782 349618 60866 349854
rect 61102 349618 96546 349854
rect 96782 349618 96866 349854
rect 97102 349618 132546 349854
rect 132782 349618 132866 349854
rect 133102 349618 168546 349854
rect 168782 349618 168866 349854
rect 169102 349618 204546 349854
rect 204782 349618 204866 349854
rect 205102 349618 240546 349854
rect 240782 349618 240866 349854
rect 241102 349618 276546 349854
rect 276782 349618 276866 349854
rect 277102 349618 312546 349854
rect 312782 349618 312866 349854
rect 313102 349618 348546 349854
rect 348782 349618 348866 349854
rect 349102 349618 384546 349854
rect 384782 349618 384866 349854
rect 385102 349618 420546 349854
rect 420782 349618 420866 349854
rect 421102 349618 456546 349854
rect 456782 349618 456866 349854
rect 457102 349618 492546 349854
rect 492782 349618 492866 349854
rect 493102 349618 528546 349854
rect 528782 349618 528866 349854
rect 529102 349618 564546 349854
rect 564782 349618 564866 349854
rect 565102 349618 591102 349854
rect 591338 349618 591422 349854
rect 591658 349618 592650 349854
rect -8726 349586 592650 349618
rect -8726 346454 592650 346486
rect -8726 346218 -6774 346454
rect -6538 346218 -6454 346454
rect -6218 346218 20826 346454
rect 21062 346218 21146 346454
rect 21382 346218 56826 346454
rect 57062 346218 57146 346454
rect 57382 346218 92826 346454
rect 93062 346218 93146 346454
rect 93382 346218 128826 346454
rect 129062 346218 129146 346454
rect 129382 346218 164826 346454
rect 165062 346218 165146 346454
rect 165382 346218 200826 346454
rect 201062 346218 201146 346454
rect 201382 346218 236826 346454
rect 237062 346218 237146 346454
rect 237382 346218 272826 346454
rect 273062 346218 273146 346454
rect 273382 346218 308826 346454
rect 309062 346218 309146 346454
rect 309382 346218 344826 346454
rect 345062 346218 345146 346454
rect 345382 346218 380826 346454
rect 381062 346218 381146 346454
rect 381382 346218 416826 346454
rect 417062 346218 417146 346454
rect 417382 346218 452826 346454
rect 453062 346218 453146 346454
rect 453382 346218 488826 346454
rect 489062 346218 489146 346454
rect 489382 346218 524826 346454
rect 525062 346218 525146 346454
rect 525382 346218 560826 346454
rect 561062 346218 561146 346454
rect 561382 346218 590142 346454
rect 590378 346218 590462 346454
rect 590698 346218 592650 346454
rect -8726 346134 592650 346218
rect -8726 345898 -6774 346134
rect -6538 345898 -6454 346134
rect -6218 345898 20826 346134
rect 21062 345898 21146 346134
rect 21382 345898 56826 346134
rect 57062 345898 57146 346134
rect 57382 345898 92826 346134
rect 93062 345898 93146 346134
rect 93382 345898 128826 346134
rect 129062 345898 129146 346134
rect 129382 345898 164826 346134
rect 165062 345898 165146 346134
rect 165382 345898 200826 346134
rect 201062 345898 201146 346134
rect 201382 345898 236826 346134
rect 237062 345898 237146 346134
rect 237382 345898 272826 346134
rect 273062 345898 273146 346134
rect 273382 345898 308826 346134
rect 309062 345898 309146 346134
rect 309382 345898 344826 346134
rect 345062 345898 345146 346134
rect 345382 345898 380826 346134
rect 381062 345898 381146 346134
rect 381382 345898 416826 346134
rect 417062 345898 417146 346134
rect 417382 345898 452826 346134
rect 453062 345898 453146 346134
rect 453382 345898 488826 346134
rect 489062 345898 489146 346134
rect 489382 345898 524826 346134
rect 525062 345898 525146 346134
rect 525382 345898 560826 346134
rect 561062 345898 561146 346134
rect 561382 345898 590142 346134
rect 590378 345898 590462 346134
rect 590698 345898 592650 346134
rect -8726 345866 592650 345898
rect -8726 342734 592650 342766
rect -8726 342498 -5814 342734
rect -5578 342498 -5494 342734
rect -5258 342498 17106 342734
rect 17342 342498 17426 342734
rect 17662 342498 53106 342734
rect 53342 342498 53426 342734
rect 53662 342498 89106 342734
rect 89342 342498 89426 342734
rect 89662 342498 125106 342734
rect 125342 342498 125426 342734
rect 125662 342498 161106 342734
rect 161342 342498 161426 342734
rect 161662 342498 197106 342734
rect 197342 342498 197426 342734
rect 197662 342498 233106 342734
rect 233342 342498 233426 342734
rect 233662 342498 269106 342734
rect 269342 342498 269426 342734
rect 269662 342498 305106 342734
rect 305342 342498 305426 342734
rect 305662 342498 341106 342734
rect 341342 342498 341426 342734
rect 341662 342498 377106 342734
rect 377342 342498 377426 342734
rect 377662 342498 413106 342734
rect 413342 342498 413426 342734
rect 413662 342498 449106 342734
rect 449342 342498 449426 342734
rect 449662 342498 485106 342734
rect 485342 342498 485426 342734
rect 485662 342498 521106 342734
rect 521342 342498 521426 342734
rect 521662 342498 557106 342734
rect 557342 342498 557426 342734
rect 557662 342498 589182 342734
rect 589418 342498 589502 342734
rect 589738 342498 592650 342734
rect -8726 342414 592650 342498
rect -8726 342178 -5814 342414
rect -5578 342178 -5494 342414
rect -5258 342178 17106 342414
rect 17342 342178 17426 342414
rect 17662 342178 53106 342414
rect 53342 342178 53426 342414
rect 53662 342178 89106 342414
rect 89342 342178 89426 342414
rect 89662 342178 125106 342414
rect 125342 342178 125426 342414
rect 125662 342178 161106 342414
rect 161342 342178 161426 342414
rect 161662 342178 197106 342414
rect 197342 342178 197426 342414
rect 197662 342178 233106 342414
rect 233342 342178 233426 342414
rect 233662 342178 269106 342414
rect 269342 342178 269426 342414
rect 269662 342178 305106 342414
rect 305342 342178 305426 342414
rect 305662 342178 341106 342414
rect 341342 342178 341426 342414
rect 341662 342178 377106 342414
rect 377342 342178 377426 342414
rect 377662 342178 413106 342414
rect 413342 342178 413426 342414
rect 413662 342178 449106 342414
rect 449342 342178 449426 342414
rect 449662 342178 485106 342414
rect 485342 342178 485426 342414
rect 485662 342178 521106 342414
rect 521342 342178 521426 342414
rect 521662 342178 557106 342414
rect 557342 342178 557426 342414
rect 557662 342178 589182 342414
rect 589418 342178 589502 342414
rect 589738 342178 592650 342414
rect -8726 342146 592650 342178
rect -8726 339014 592650 339046
rect -8726 338778 -4854 339014
rect -4618 338778 -4534 339014
rect -4298 338778 13386 339014
rect 13622 338778 13706 339014
rect 13942 338778 49386 339014
rect 49622 338778 49706 339014
rect 49942 338778 85386 339014
rect 85622 338778 85706 339014
rect 85942 338778 121386 339014
rect 121622 338778 121706 339014
rect 121942 338778 157386 339014
rect 157622 338778 157706 339014
rect 157942 338778 193386 339014
rect 193622 338778 193706 339014
rect 193942 338778 229386 339014
rect 229622 338778 229706 339014
rect 229942 338778 265386 339014
rect 265622 338778 265706 339014
rect 265942 338778 301386 339014
rect 301622 338778 301706 339014
rect 301942 338778 337386 339014
rect 337622 338778 337706 339014
rect 337942 338778 373386 339014
rect 373622 338778 373706 339014
rect 373942 338778 409386 339014
rect 409622 338778 409706 339014
rect 409942 338778 445386 339014
rect 445622 338778 445706 339014
rect 445942 338778 481386 339014
rect 481622 338778 481706 339014
rect 481942 338778 517386 339014
rect 517622 338778 517706 339014
rect 517942 338778 553386 339014
rect 553622 338778 553706 339014
rect 553942 338778 588222 339014
rect 588458 338778 588542 339014
rect 588778 338778 592650 339014
rect -8726 338694 592650 338778
rect -8726 338458 -4854 338694
rect -4618 338458 -4534 338694
rect -4298 338458 13386 338694
rect 13622 338458 13706 338694
rect 13942 338458 49386 338694
rect 49622 338458 49706 338694
rect 49942 338458 85386 338694
rect 85622 338458 85706 338694
rect 85942 338458 121386 338694
rect 121622 338458 121706 338694
rect 121942 338458 157386 338694
rect 157622 338458 157706 338694
rect 157942 338458 193386 338694
rect 193622 338458 193706 338694
rect 193942 338458 229386 338694
rect 229622 338458 229706 338694
rect 229942 338458 265386 338694
rect 265622 338458 265706 338694
rect 265942 338458 301386 338694
rect 301622 338458 301706 338694
rect 301942 338458 337386 338694
rect 337622 338458 337706 338694
rect 337942 338458 373386 338694
rect 373622 338458 373706 338694
rect 373942 338458 409386 338694
rect 409622 338458 409706 338694
rect 409942 338458 445386 338694
rect 445622 338458 445706 338694
rect 445942 338458 481386 338694
rect 481622 338458 481706 338694
rect 481942 338458 517386 338694
rect 517622 338458 517706 338694
rect 517942 338458 553386 338694
rect 553622 338458 553706 338694
rect 553942 338458 588222 338694
rect 588458 338458 588542 338694
rect 588778 338458 592650 338694
rect -8726 338426 592650 338458
rect -8726 335294 592650 335326
rect -8726 335058 -3894 335294
rect -3658 335058 -3574 335294
rect -3338 335058 9666 335294
rect 9902 335058 9986 335294
rect 10222 335058 45666 335294
rect 45902 335058 45986 335294
rect 46222 335058 81666 335294
rect 81902 335058 81986 335294
rect 82222 335058 117666 335294
rect 117902 335058 117986 335294
rect 118222 335058 153666 335294
rect 153902 335058 153986 335294
rect 154222 335058 189666 335294
rect 189902 335058 189986 335294
rect 190222 335058 225666 335294
rect 225902 335058 225986 335294
rect 226222 335058 261666 335294
rect 261902 335058 261986 335294
rect 262222 335058 297666 335294
rect 297902 335058 297986 335294
rect 298222 335058 333666 335294
rect 333902 335058 333986 335294
rect 334222 335058 369666 335294
rect 369902 335058 369986 335294
rect 370222 335058 405666 335294
rect 405902 335058 405986 335294
rect 406222 335058 441666 335294
rect 441902 335058 441986 335294
rect 442222 335058 477666 335294
rect 477902 335058 477986 335294
rect 478222 335058 513666 335294
rect 513902 335058 513986 335294
rect 514222 335058 549666 335294
rect 549902 335058 549986 335294
rect 550222 335058 587262 335294
rect 587498 335058 587582 335294
rect 587818 335058 592650 335294
rect -8726 334974 592650 335058
rect -8726 334738 -3894 334974
rect -3658 334738 -3574 334974
rect -3338 334738 9666 334974
rect 9902 334738 9986 334974
rect 10222 334738 45666 334974
rect 45902 334738 45986 334974
rect 46222 334738 81666 334974
rect 81902 334738 81986 334974
rect 82222 334738 117666 334974
rect 117902 334738 117986 334974
rect 118222 334738 153666 334974
rect 153902 334738 153986 334974
rect 154222 334738 189666 334974
rect 189902 334738 189986 334974
rect 190222 334738 225666 334974
rect 225902 334738 225986 334974
rect 226222 334738 261666 334974
rect 261902 334738 261986 334974
rect 262222 334738 297666 334974
rect 297902 334738 297986 334974
rect 298222 334738 333666 334974
rect 333902 334738 333986 334974
rect 334222 334738 369666 334974
rect 369902 334738 369986 334974
rect 370222 334738 405666 334974
rect 405902 334738 405986 334974
rect 406222 334738 441666 334974
rect 441902 334738 441986 334974
rect 442222 334738 477666 334974
rect 477902 334738 477986 334974
rect 478222 334738 513666 334974
rect 513902 334738 513986 334974
rect 514222 334738 549666 334974
rect 549902 334738 549986 334974
rect 550222 334738 587262 334974
rect 587498 334738 587582 334974
rect 587818 334738 592650 334974
rect -8726 334706 592650 334738
rect -8726 331574 592650 331606
rect -8726 331338 -2934 331574
rect -2698 331338 -2614 331574
rect -2378 331338 5946 331574
rect 6182 331338 6266 331574
rect 6502 331338 41946 331574
rect 42182 331338 42266 331574
rect 42502 331338 77946 331574
rect 78182 331338 78266 331574
rect 78502 331338 113946 331574
rect 114182 331338 114266 331574
rect 114502 331338 149946 331574
rect 150182 331338 150266 331574
rect 150502 331338 185946 331574
rect 186182 331338 186266 331574
rect 186502 331338 221946 331574
rect 222182 331338 222266 331574
rect 222502 331338 257946 331574
rect 258182 331338 258266 331574
rect 258502 331338 293946 331574
rect 294182 331338 294266 331574
rect 294502 331338 329946 331574
rect 330182 331338 330266 331574
rect 330502 331338 365946 331574
rect 366182 331338 366266 331574
rect 366502 331338 401946 331574
rect 402182 331338 402266 331574
rect 402502 331338 437946 331574
rect 438182 331338 438266 331574
rect 438502 331338 473946 331574
rect 474182 331338 474266 331574
rect 474502 331338 509946 331574
rect 510182 331338 510266 331574
rect 510502 331338 545946 331574
rect 546182 331338 546266 331574
rect 546502 331338 581946 331574
rect 582182 331338 582266 331574
rect 582502 331338 586302 331574
rect 586538 331338 586622 331574
rect 586858 331338 592650 331574
rect -8726 331254 592650 331338
rect -8726 331018 -2934 331254
rect -2698 331018 -2614 331254
rect -2378 331018 5946 331254
rect 6182 331018 6266 331254
rect 6502 331018 41946 331254
rect 42182 331018 42266 331254
rect 42502 331018 77946 331254
rect 78182 331018 78266 331254
rect 78502 331018 113946 331254
rect 114182 331018 114266 331254
rect 114502 331018 149946 331254
rect 150182 331018 150266 331254
rect 150502 331018 185946 331254
rect 186182 331018 186266 331254
rect 186502 331018 221946 331254
rect 222182 331018 222266 331254
rect 222502 331018 257946 331254
rect 258182 331018 258266 331254
rect 258502 331018 293946 331254
rect 294182 331018 294266 331254
rect 294502 331018 329946 331254
rect 330182 331018 330266 331254
rect 330502 331018 365946 331254
rect 366182 331018 366266 331254
rect 366502 331018 401946 331254
rect 402182 331018 402266 331254
rect 402502 331018 437946 331254
rect 438182 331018 438266 331254
rect 438502 331018 473946 331254
rect 474182 331018 474266 331254
rect 474502 331018 509946 331254
rect 510182 331018 510266 331254
rect 510502 331018 545946 331254
rect 546182 331018 546266 331254
rect 546502 331018 581946 331254
rect 582182 331018 582266 331254
rect 582502 331018 586302 331254
rect 586538 331018 586622 331254
rect 586858 331018 592650 331254
rect -8726 330986 592650 331018
rect -8726 327854 592650 327886
rect -8726 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 2226 327854
rect 2462 327618 2546 327854
rect 2782 327618 38226 327854
rect 38462 327618 38546 327854
rect 38782 327618 74226 327854
rect 74462 327618 74546 327854
rect 74782 327618 110226 327854
rect 110462 327618 110546 327854
rect 110782 327618 146226 327854
rect 146462 327618 146546 327854
rect 146782 327618 182226 327854
rect 182462 327618 182546 327854
rect 182782 327618 218226 327854
rect 218462 327618 218546 327854
rect 218782 327618 254226 327854
rect 254462 327618 254546 327854
rect 254782 327618 290226 327854
rect 290462 327618 290546 327854
rect 290782 327618 326226 327854
rect 326462 327618 326546 327854
rect 326782 327618 362226 327854
rect 362462 327618 362546 327854
rect 362782 327618 398226 327854
rect 398462 327618 398546 327854
rect 398782 327618 434226 327854
rect 434462 327618 434546 327854
rect 434782 327618 470226 327854
rect 470462 327618 470546 327854
rect 470782 327618 506226 327854
rect 506462 327618 506546 327854
rect 506782 327618 542226 327854
rect 542462 327618 542546 327854
rect 542782 327618 578226 327854
rect 578462 327618 578546 327854
rect 578782 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 592650 327854
rect -8726 327534 592650 327618
rect -8726 327298 -1974 327534
rect -1738 327298 -1654 327534
rect -1418 327298 2226 327534
rect 2462 327298 2546 327534
rect 2782 327298 38226 327534
rect 38462 327298 38546 327534
rect 38782 327298 74226 327534
rect 74462 327298 74546 327534
rect 74782 327298 110226 327534
rect 110462 327298 110546 327534
rect 110782 327298 146226 327534
rect 146462 327298 146546 327534
rect 146782 327298 182226 327534
rect 182462 327298 182546 327534
rect 182782 327298 218226 327534
rect 218462 327298 218546 327534
rect 218782 327298 254226 327534
rect 254462 327298 254546 327534
rect 254782 327298 290226 327534
rect 290462 327298 290546 327534
rect 290782 327298 326226 327534
rect 326462 327298 326546 327534
rect 326782 327298 362226 327534
rect 362462 327298 362546 327534
rect 362782 327298 398226 327534
rect 398462 327298 398546 327534
rect 398782 327298 434226 327534
rect 434462 327298 434546 327534
rect 434782 327298 470226 327534
rect 470462 327298 470546 327534
rect 470782 327298 506226 327534
rect 506462 327298 506546 327534
rect 506782 327298 542226 327534
rect 542462 327298 542546 327534
rect 542782 327298 578226 327534
rect 578462 327298 578546 327534
rect 578782 327298 585342 327534
rect 585578 327298 585662 327534
rect 585898 327298 592650 327534
rect -8726 327266 592650 327298
rect -8726 317894 592650 317926
rect -8726 317658 -8694 317894
rect -8458 317658 -8374 317894
rect -8138 317658 28266 317894
rect 28502 317658 28586 317894
rect 28822 317658 64266 317894
rect 64502 317658 64586 317894
rect 64822 317658 100266 317894
rect 100502 317658 100586 317894
rect 100822 317658 136266 317894
rect 136502 317658 136586 317894
rect 136822 317658 172266 317894
rect 172502 317658 172586 317894
rect 172822 317658 208266 317894
rect 208502 317658 208586 317894
rect 208822 317658 244266 317894
rect 244502 317658 244586 317894
rect 244822 317658 280266 317894
rect 280502 317658 280586 317894
rect 280822 317658 316266 317894
rect 316502 317658 316586 317894
rect 316822 317658 352266 317894
rect 352502 317658 352586 317894
rect 352822 317658 388266 317894
rect 388502 317658 388586 317894
rect 388822 317658 424266 317894
rect 424502 317658 424586 317894
rect 424822 317658 460266 317894
rect 460502 317658 460586 317894
rect 460822 317658 496266 317894
rect 496502 317658 496586 317894
rect 496822 317658 532266 317894
rect 532502 317658 532586 317894
rect 532822 317658 568266 317894
rect 568502 317658 568586 317894
rect 568822 317658 592062 317894
rect 592298 317658 592382 317894
rect 592618 317658 592650 317894
rect -8726 317574 592650 317658
rect -8726 317338 -8694 317574
rect -8458 317338 -8374 317574
rect -8138 317338 28266 317574
rect 28502 317338 28586 317574
rect 28822 317338 64266 317574
rect 64502 317338 64586 317574
rect 64822 317338 100266 317574
rect 100502 317338 100586 317574
rect 100822 317338 136266 317574
rect 136502 317338 136586 317574
rect 136822 317338 172266 317574
rect 172502 317338 172586 317574
rect 172822 317338 208266 317574
rect 208502 317338 208586 317574
rect 208822 317338 244266 317574
rect 244502 317338 244586 317574
rect 244822 317338 280266 317574
rect 280502 317338 280586 317574
rect 280822 317338 316266 317574
rect 316502 317338 316586 317574
rect 316822 317338 352266 317574
rect 352502 317338 352586 317574
rect 352822 317338 388266 317574
rect 388502 317338 388586 317574
rect 388822 317338 424266 317574
rect 424502 317338 424586 317574
rect 424822 317338 460266 317574
rect 460502 317338 460586 317574
rect 460822 317338 496266 317574
rect 496502 317338 496586 317574
rect 496822 317338 532266 317574
rect 532502 317338 532586 317574
rect 532822 317338 568266 317574
rect 568502 317338 568586 317574
rect 568822 317338 592062 317574
rect 592298 317338 592382 317574
rect 592618 317338 592650 317574
rect -8726 317306 592650 317338
rect -8726 314174 592650 314206
rect -8726 313938 -7734 314174
rect -7498 313938 -7414 314174
rect -7178 313938 24546 314174
rect 24782 313938 24866 314174
rect 25102 313938 60546 314174
rect 60782 313938 60866 314174
rect 61102 313938 96546 314174
rect 96782 313938 96866 314174
rect 97102 313938 132546 314174
rect 132782 313938 132866 314174
rect 133102 313938 168546 314174
rect 168782 313938 168866 314174
rect 169102 313938 204546 314174
rect 204782 313938 204866 314174
rect 205102 313938 240546 314174
rect 240782 313938 240866 314174
rect 241102 313938 276546 314174
rect 276782 313938 276866 314174
rect 277102 313938 312546 314174
rect 312782 313938 312866 314174
rect 313102 313938 348546 314174
rect 348782 313938 348866 314174
rect 349102 313938 384546 314174
rect 384782 313938 384866 314174
rect 385102 313938 420546 314174
rect 420782 313938 420866 314174
rect 421102 313938 456546 314174
rect 456782 313938 456866 314174
rect 457102 313938 492546 314174
rect 492782 313938 492866 314174
rect 493102 313938 528546 314174
rect 528782 313938 528866 314174
rect 529102 313938 564546 314174
rect 564782 313938 564866 314174
rect 565102 313938 591102 314174
rect 591338 313938 591422 314174
rect 591658 313938 592650 314174
rect -8726 313854 592650 313938
rect -8726 313618 -7734 313854
rect -7498 313618 -7414 313854
rect -7178 313618 24546 313854
rect 24782 313618 24866 313854
rect 25102 313618 60546 313854
rect 60782 313618 60866 313854
rect 61102 313618 96546 313854
rect 96782 313618 96866 313854
rect 97102 313618 132546 313854
rect 132782 313618 132866 313854
rect 133102 313618 168546 313854
rect 168782 313618 168866 313854
rect 169102 313618 204546 313854
rect 204782 313618 204866 313854
rect 205102 313618 240546 313854
rect 240782 313618 240866 313854
rect 241102 313618 276546 313854
rect 276782 313618 276866 313854
rect 277102 313618 312546 313854
rect 312782 313618 312866 313854
rect 313102 313618 348546 313854
rect 348782 313618 348866 313854
rect 349102 313618 384546 313854
rect 384782 313618 384866 313854
rect 385102 313618 420546 313854
rect 420782 313618 420866 313854
rect 421102 313618 456546 313854
rect 456782 313618 456866 313854
rect 457102 313618 492546 313854
rect 492782 313618 492866 313854
rect 493102 313618 528546 313854
rect 528782 313618 528866 313854
rect 529102 313618 564546 313854
rect 564782 313618 564866 313854
rect 565102 313618 591102 313854
rect 591338 313618 591422 313854
rect 591658 313618 592650 313854
rect -8726 313586 592650 313618
rect -8726 310454 592650 310486
rect -8726 310218 -6774 310454
rect -6538 310218 -6454 310454
rect -6218 310218 20826 310454
rect 21062 310218 21146 310454
rect 21382 310218 56826 310454
rect 57062 310218 57146 310454
rect 57382 310218 92826 310454
rect 93062 310218 93146 310454
rect 93382 310218 128826 310454
rect 129062 310218 129146 310454
rect 129382 310218 164826 310454
rect 165062 310218 165146 310454
rect 165382 310218 200826 310454
rect 201062 310218 201146 310454
rect 201382 310218 236826 310454
rect 237062 310218 237146 310454
rect 237382 310218 272826 310454
rect 273062 310218 273146 310454
rect 273382 310218 308826 310454
rect 309062 310218 309146 310454
rect 309382 310218 344826 310454
rect 345062 310218 345146 310454
rect 345382 310218 380826 310454
rect 381062 310218 381146 310454
rect 381382 310218 416826 310454
rect 417062 310218 417146 310454
rect 417382 310218 452826 310454
rect 453062 310218 453146 310454
rect 453382 310218 488826 310454
rect 489062 310218 489146 310454
rect 489382 310218 524826 310454
rect 525062 310218 525146 310454
rect 525382 310218 560826 310454
rect 561062 310218 561146 310454
rect 561382 310218 590142 310454
rect 590378 310218 590462 310454
rect 590698 310218 592650 310454
rect -8726 310134 592650 310218
rect -8726 309898 -6774 310134
rect -6538 309898 -6454 310134
rect -6218 309898 20826 310134
rect 21062 309898 21146 310134
rect 21382 309898 56826 310134
rect 57062 309898 57146 310134
rect 57382 309898 92826 310134
rect 93062 309898 93146 310134
rect 93382 309898 128826 310134
rect 129062 309898 129146 310134
rect 129382 309898 164826 310134
rect 165062 309898 165146 310134
rect 165382 309898 200826 310134
rect 201062 309898 201146 310134
rect 201382 309898 236826 310134
rect 237062 309898 237146 310134
rect 237382 309898 272826 310134
rect 273062 309898 273146 310134
rect 273382 309898 308826 310134
rect 309062 309898 309146 310134
rect 309382 309898 344826 310134
rect 345062 309898 345146 310134
rect 345382 309898 380826 310134
rect 381062 309898 381146 310134
rect 381382 309898 416826 310134
rect 417062 309898 417146 310134
rect 417382 309898 452826 310134
rect 453062 309898 453146 310134
rect 453382 309898 488826 310134
rect 489062 309898 489146 310134
rect 489382 309898 524826 310134
rect 525062 309898 525146 310134
rect 525382 309898 560826 310134
rect 561062 309898 561146 310134
rect 561382 309898 590142 310134
rect 590378 309898 590462 310134
rect 590698 309898 592650 310134
rect -8726 309866 592650 309898
rect -8726 306734 592650 306766
rect -8726 306498 -5814 306734
rect -5578 306498 -5494 306734
rect -5258 306498 17106 306734
rect 17342 306498 17426 306734
rect 17662 306498 53106 306734
rect 53342 306498 53426 306734
rect 53662 306498 89106 306734
rect 89342 306498 89426 306734
rect 89662 306498 125106 306734
rect 125342 306498 125426 306734
rect 125662 306498 161106 306734
rect 161342 306498 161426 306734
rect 161662 306498 197106 306734
rect 197342 306498 197426 306734
rect 197662 306498 233106 306734
rect 233342 306498 233426 306734
rect 233662 306498 269106 306734
rect 269342 306498 269426 306734
rect 269662 306498 305106 306734
rect 305342 306498 305426 306734
rect 305662 306498 341106 306734
rect 341342 306498 341426 306734
rect 341662 306498 377106 306734
rect 377342 306498 377426 306734
rect 377662 306498 413106 306734
rect 413342 306498 413426 306734
rect 413662 306498 449106 306734
rect 449342 306498 449426 306734
rect 449662 306498 485106 306734
rect 485342 306498 485426 306734
rect 485662 306498 521106 306734
rect 521342 306498 521426 306734
rect 521662 306498 557106 306734
rect 557342 306498 557426 306734
rect 557662 306498 589182 306734
rect 589418 306498 589502 306734
rect 589738 306498 592650 306734
rect -8726 306414 592650 306498
rect -8726 306178 -5814 306414
rect -5578 306178 -5494 306414
rect -5258 306178 17106 306414
rect 17342 306178 17426 306414
rect 17662 306178 53106 306414
rect 53342 306178 53426 306414
rect 53662 306178 89106 306414
rect 89342 306178 89426 306414
rect 89662 306178 125106 306414
rect 125342 306178 125426 306414
rect 125662 306178 161106 306414
rect 161342 306178 161426 306414
rect 161662 306178 197106 306414
rect 197342 306178 197426 306414
rect 197662 306178 233106 306414
rect 233342 306178 233426 306414
rect 233662 306178 269106 306414
rect 269342 306178 269426 306414
rect 269662 306178 305106 306414
rect 305342 306178 305426 306414
rect 305662 306178 341106 306414
rect 341342 306178 341426 306414
rect 341662 306178 377106 306414
rect 377342 306178 377426 306414
rect 377662 306178 413106 306414
rect 413342 306178 413426 306414
rect 413662 306178 449106 306414
rect 449342 306178 449426 306414
rect 449662 306178 485106 306414
rect 485342 306178 485426 306414
rect 485662 306178 521106 306414
rect 521342 306178 521426 306414
rect 521662 306178 557106 306414
rect 557342 306178 557426 306414
rect 557662 306178 589182 306414
rect 589418 306178 589502 306414
rect 589738 306178 592650 306414
rect -8726 306146 592650 306178
rect -8726 303014 592650 303046
rect -8726 302778 -4854 303014
rect -4618 302778 -4534 303014
rect -4298 302778 13386 303014
rect 13622 302778 13706 303014
rect 13942 302778 49386 303014
rect 49622 302778 49706 303014
rect 49942 302778 85386 303014
rect 85622 302778 85706 303014
rect 85942 302778 121386 303014
rect 121622 302778 121706 303014
rect 121942 302778 157386 303014
rect 157622 302778 157706 303014
rect 157942 302778 193386 303014
rect 193622 302778 193706 303014
rect 193942 302778 229386 303014
rect 229622 302778 229706 303014
rect 229942 302778 265386 303014
rect 265622 302778 265706 303014
rect 265942 302778 301386 303014
rect 301622 302778 301706 303014
rect 301942 302778 337386 303014
rect 337622 302778 337706 303014
rect 337942 302778 373386 303014
rect 373622 302778 373706 303014
rect 373942 302778 409386 303014
rect 409622 302778 409706 303014
rect 409942 302778 445386 303014
rect 445622 302778 445706 303014
rect 445942 302778 481386 303014
rect 481622 302778 481706 303014
rect 481942 302778 517386 303014
rect 517622 302778 517706 303014
rect 517942 302778 553386 303014
rect 553622 302778 553706 303014
rect 553942 302778 588222 303014
rect 588458 302778 588542 303014
rect 588778 302778 592650 303014
rect -8726 302694 592650 302778
rect -8726 302458 -4854 302694
rect -4618 302458 -4534 302694
rect -4298 302458 13386 302694
rect 13622 302458 13706 302694
rect 13942 302458 49386 302694
rect 49622 302458 49706 302694
rect 49942 302458 85386 302694
rect 85622 302458 85706 302694
rect 85942 302458 121386 302694
rect 121622 302458 121706 302694
rect 121942 302458 157386 302694
rect 157622 302458 157706 302694
rect 157942 302458 193386 302694
rect 193622 302458 193706 302694
rect 193942 302458 229386 302694
rect 229622 302458 229706 302694
rect 229942 302458 265386 302694
rect 265622 302458 265706 302694
rect 265942 302458 301386 302694
rect 301622 302458 301706 302694
rect 301942 302458 337386 302694
rect 337622 302458 337706 302694
rect 337942 302458 373386 302694
rect 373622 302458 373706 302694
rect 373942 302458 409386 302694
rect 409622 302458 409706 302694
rect 409942 302458 445386 302694
rect 445622 302458 445706 302694
rect 445942 302458 481386 302694
rect 481622 302458 481706 302694
rect 481942 302458 517386 302694
rect 517622 302458 517706 302694
rect 517942 302458 553386 302694
rect 553622 302458 553706 302694
rect 553942 302458 588222 302694
rect 588458 302458 588542 302694
rect 588778 302458 592650 302694
rect -8726 302426 592650 302458
rect -8726 299294 592650 299326
rect -8726 299058 -3894 299294
rect -3658 299058 -3574 299294
rect -3338 299058 9666 299294
rect 9902 299058 9986 299294
rect 10222 299058 45666 299294
rect 45902 299058 45986 299294
rect 46222 299058 81666 299294
rect 81902 299058 81986 299294
rect 82222 299058 117666 299294
rect 117902 299058 117986 299294
rect 118222 299058 153666 299294
rect 153902 299058 153986 299294
rect 154222 299058 189666 299294
rect 189902 299058 189986 299294
rect 190222 299058 225666 299294
rect 225902 299058 225986 299294
rect 226222 299058 261666 299294
rect 261902 299058 261986 299294
rect 262222 299058 297666 299294
rect 297902 299058 297986 299294
rect 298222 299058 333666 299294
rect 333902 299058 333986 299294
rect 334222 299058 369666 299294
rect 369902 299058 369986 299294
rect 370222 299058 405666 299294
rect 405902 299058 405986 299294
rect 406222 299058 441666 299294
rect 441902 299058 441986 299294
rect 442222 299058 477666 299294
rect 477902 299058 477986 299294
rect 478222 299058 513666 299294
rect 513902 299058 513986 299294
rect 514222 299058 549666 299294
rect 549902 299058 549986 299294
rect 550222 299058 587262 299294
rect 587498 299058 587582 299294
rect 587818 299058 592650 299294
rect -8726 298974 592650 299058
rect -8726 298738 -3894 298974
rect -3658 298738 -3574 298974
rect -3338 298738 9666 298974
rect 9902 298738 9986 298974
rect 10222 298738 45666 298974
rect 45902 298738 45986 298974
rect 46222 298738 81666 298974
rect 81902 298738 81986 298974
rect 82222 298738 117666 298974
rect 117902 298738 117986 298974
rect 118222 298738 153666 298974
rect 153902 298738 153986 298974
rect 154222 298738 189666 298974
rect 189902 298738 189986 298974
rect 190222 298738 225666 298974
rect 225902 298738 225986 298974
rect 226222 298738 261666 298974
rect 261902 298738 261986 298974
rect 262222 298738 297666 298974
rect 297902 298738 297986 298974
rect 298222 298738 333666 298974
rect 333902 298738 333986 298974
rect 334222 298738 369666 298974
rect 369902 298738 369986 298974
rect 370222 298738 405666 298974
rect 405902 298738 405986 298974
rect 406222 298738 441666 298974
rect 441902 298738 441986 298974
rect 442222 298738 477666 298974
rect 477902 298738 477986 298974
rect 478222 298738 513666 298974
rect 513902 298738 513986 298974
rect 514222 298738 549666 298974
rect 549902 298738 549986 298974
rect 550222 298738 587262 298974
rect 587498 298738 587582 298974
rect 587818 298738 592650 298974
rect -8726 298706 592650 298738
rect -8726 295574 592650 295606
rect -8726 295338 -2934 295574
rect -2698 295338 -2614 295574
rect -2378 295338 5946 295574
rect 6182 295338 6266 295574
rect 6502 295338 41946 295574
rect 42182 295338 42266 295574
rect 42502 295338 77946 295574
rect 78182 295338 78266 295574
rect 78502 295338 113946 295574
rect 114182 295338 114266 295574
rect 114502 295338 149946 295574
rect 150182 295338 150266 295574
rect 150502 295338 185946 295574
rect 186182 295338 186266 295574
rect 186502 295338 221946 295574
rect 222182 295338 222266 295574
rect 222502 295338 257946 295574
rect 258182 295338 258266 295574
rect 258502 295338 293946 295574
rect 294182 295338 294266 295574
rect 294502 295338 329946 295574
rect 330182 295338 330266 295574
rect 330502 295338 365946 295574
rect 366182 295338 366266 295574
rect 366502 295338 401946 295574
rect 402182 295338 402266 295574
rect 402502 295338 437946 295574
rect 438182 295338 438266 295574
rect 438502 295338 473946 295574
rect 474182 295338 474266 295574
rect 474502 295338 509946 295574
rect 510182 295338 510266 295574
rect 510502 295338 545946 295574
rect 546182 295338 546266 295574
rect 546502 295338 581946 295574
rect 582182 295338 582266 295574
rect 582502 295338 586302 295574
rect 586538 295338 586622 295574
rect 586858 295338 592650 295574
rect -8726 295254 592650 295338
rect -8726 295018 -2934 295254
rect -2698 295018 -2614 295254
rect -2378 295018 5946 295254
rect 6182 295018 6266 295254
rect 6502 295018 41946 295254
rect 42182 295018 42266 295254
rect 42502 295018 77946 295254
rect 78182 295018 78266 295254
rect 78502 295018 113946 295254
rect 114182 295018 114266 295254
rect 114502 295018 149946 295254
rect 150182 295018 150266 295254
rect 150502 295018 185946 295254
rect 186182 295018 186266 295254
rect 186502 295018 221946 295254
rect 222182 295018 222266 295254
rect 222502 295018 257946 295254
rect 258182 295018 258266 295254
rect 258502 295018 293946 295254
rect 294182 295018 294266 295254
rect 294502 295018 329946 295254
rect 330182 295018 330266 295254
rect 330502 295018 365946 295254
rect 366182 295018 366266 295254
rect 366502 295018 401946 295254
rect 402182 295018 402266 295254
rect 402502 295018 437946 295254
rect 438182 295018 438266 295254
rect 438502 295018 473946 295254
rect 474182 295018 474266 295254
rect 474502 295018 509946 295254
rect 510182 295018 510266 295254
rect 510502 295018 545946 295254
rect 546182 295018 546266 295254
rect 546502 295018 581946 295254
rect 582182 295018 582266 295254
rect 582502 295018 586302 295254
rect 586538 295018 586622 295254
rect 586858 295018 592650 295254
rect -8726 294986 592650 295018
rect -8726 291854 592650 291886
rect -8726 291618 -1974 291854
rect -1738 291618 -1654 291854
rect -1418 291618 2226 291854
rect 2462 291618 2546 291854
rect 2782 291618 38226 291854
rect 38462 291618 38546 291854
rect 38782 291618 74226 291854
rect 74462 291618 74546 291854
rect 74782 291618 110226 291854
rect 110462 291618 110546 291854
rect 110782 291618 146226 291854
rect 146462 291618 146546 291854
rect 146782 291618 182226 291854
rect 182462 291618 182546 291854
rect 182782 291618 218226 291854
rect 218462 291618 218546 291854
rect 218782 291618 254226 291854
rect 254462 291618 254546 291854
rect 254782 291618 290226 291854
rect 290462 291618 290546 291854
rect 290782 291618 326226 291854
rect 326462 291618 326546 291854
rect 326782 291618 362226 291854
rect 362462 291618 362546 291854
rect 362782 291618 398226 291854
rect 398462 291618 398546 291854
rect 398782 291618 434226 291854
rect 434462 291618 434546 291854
rect 434782 291618 470226 291854
rect 470462 291618 470546 291854
rect 470782 291618 506226 291854
rect 506462 291618 506546 291854
rect 506782 291618 542226 291854
rect 542462 291618 542546 291854
rect 542782 291618 578226 291854
rect 578462 291618 578546 291854
rect 578782 291618 585342 291854
rect 585578 291618 585662 291854
rect 585898 291618 592650 291854
rect -8726 291534 592650 291618
rect -8726 291298 -1974 291534
rect -1738 291298 -1654 291534
rect -1418 291298 2226 291534
rect 2462 291298 2546 291534
rect 2782 291298 38226 291534
rect 38462 291298 38546 291534
rect 38782 291298 74226 291534
rect 74462 291298 74546 291534
rect 74782 291298 110226 291534
rect 110462 291298 110546 291534
rect 110782 291298 146226 291534
rect 146462 291298 146546 291534
rect 146782 291298 182226 291534
rect 182462 291298 182546 291534
rect 182782 291298 218226 291534
rect 218462 291298 218546 291534
rect 218782 291298 254226 291534
rect 254462 291298 254546 291534
rect 254782 291298 290226 291534
rect 290462 291298 290546 291534
rect 290782 291298 326226 291534
rect 326462 291298 326546 291534
rect 326782 291298 362226 291534
rect 362462 291298 362546 291534
rect 362782 291298 398226 291534
rect 398462 291298 398546 291534
rect 398782 291298 434226 291534
rect 434462 291298 434546 291534
rect 434782 291298 470226 291534
rect 470462 291298 470546 291534
rect 470782 291298 506226 291534
rect 506462 291298 506546 291534
rect 506782 291298 542226 291534
rect 542462 291298 542546 291534
rect 542782 291298 578226 291534
rect 578462 291298 578546 291534
rect 578782 291298 585342 291534
rect 585578 291298 585662 291534
rect 585898 291298 592650 291534
rect -8726 291266 592650 291298
rect -8726 281894 592650 281926
rect -8726 281658 -8694 281894
rect -8458 281658 -8374 281894
rect -8138 281658 28266 281894
rect 28502 281658 28586 281894
rect 28822 281658 64266 281894
rect 64502 281658 64586 281894
rect 64822 281658 100266 281894
rect 100502 281658 100586 281894
rect 100822 281658 136266 281894
rect 136502 281658 136586 281894
rect 136822 281658 172266 281894
rect 172502 281658 172586 281894
rect 172822 281658 208266 281894
rect 208502 281658 208586 281894
rect 208822 281658 244266 281894
rect 244502 281658 244586 281894
rect 244822 281658 280266 281894
rect 280502 281658 280586 281894
rect 280822 281658 316266 281894
rect 316502 281658 316586 281894
rect 316822 281658 352266 281894
rect 352502 281658 352586 281894
rect 352822 281658 388266 281894
rect 388502 281658 388586 281894
rect 388822 281658 424266 281894
rect 424502 281658 424586 281894
rect 424822 281658 460266 281894
rect 460502 281658 460586 281894
rect 460822 281658 496266 281894
rect 496502 281658 496586 281894
rect 496822 281658 532266 281894
rect 532502 281658 532586 281894
rect 532822 281658 568266 281894
rect 568502 281658 568586 281894
rect 568822 281658 592062 281894
rect 592298 281658 592382 281894
rect 592618 281658 592650 281894
rect -8726 281574 592650 281658
rect -8726 281338 -8694 281574
rect -8458 281338 -8374 281574
rect -8138 281338 28266 281574
rect 28502 281338 28586 281574
rect 28822 281338 64266 281574
rect 64502 281338 64586 281574
rect 64822 281338 100266 281574
rect 100502 281338 100586 281574
rect 100822 281338 136266 281574
rect 136502 281338 136586 281574
rect 136822 281338 172266 281574
rect 172502 281338 172586 281574
rect 172822 281338 208266 281574
rect 208502 281338 208586 281574
rect 208822 281338 244266 281574
rect 244502 281338 244586 281574
rect 244822 281338 280266 281574
rect 280502 281338 280586 281574
rect 280822 281338 316266 281574
rect 316502 281338 316586 281574
rect 316822 281338 352266 281574
rect 352502 281338 352586 281574
rect 352822 281338 388266 281574
rect 388502 281338 388586 281574
rect 388822 281338 424266 281574
rect 424502 281338 424586 281574
rect 424822 281338 460266 281574
rect 460502 281338 460586 281574
rect 460822 281338 496266 281574
rect 496502 281338 496586 281574
rect 496822 281338 532266 281574
rect 532502 281338 532586 281574
rect 532822 281338 568266 281574
rect 568502 281338 568586 281574
rect 568822 281338 592062 281574
rect 592298 281338 592382 281574
rect 592618 281338 592650 281574
rect -8726 281306 592650 281338
rect -8726 278174 592650 278206
rect -8726 277938 -7734 278174
rect -7498 277938 -7414 278174
rect -7178 277938 24546 278174
rect 24782 277938 24866 278174
rect 25102 277938 60546 278174
rect 60782 277938 60866 278174
rect 61102 277938 96546 278174
rect 96782 277938 96866 278174
rect 97102 277938 132546 278174
rect 132782 277938 132866 278174
rect 133102 277938 168546 278174
rect 168782 277938 168866 278174
rect 169102 277938 204546 278174
rect 204782 277938 204866 278174
rect 205102 277938 240546 278174
rect 240782 277938 240866 278174
rect 241102 277938 276546 278174
rect 276782 277938 276866 278174
rect 277102 277938 312546 278174
rect 312782 277938 312866 278174
rect 313102 277938 348546 278174
rect 348782 277938 348866 278174
rect 349102 277938 384546 278174
rect 384782 277938 384866 278174
rect 385102 277938 420546 278174
rect 420782 277938 420866 278174
rect 421102 277938 456546 278174
rect 456782 277938 456866 278174
rect 457102 277938 492546 278174
rect 492782 277938 492866 278174
rect 493102 277938 528546 278174
rect 528782 277938 528866 278174
rect 529102 277938 564546 278174
rect 564782 277938 564866 278174
rect 565102 277938 591102 278174
rect 591338 277938 591422 278174
rect 591658 277938 592650 278174
rect -8726 277854 592650 277938
rect -8726 277618 -7734 277854
rect -7498 277618 -7414 277854
rect -7178 277618 24546 277854
rect 24782 277618 24866 277854
rect 25102 277618 60546 277854
rect 60782 277618 60866 277854
rect 61102 277618 96546 277854
rect 96782 277618 96866 277854
rect 97102 277618 132546 277854
rect 132782 277618 132866 277854
rect 133102 277618 168546 277854
rect 168782 277618 168866 277854
rect 169102 277618 204546 277854
rect 204782 277618 204866 277854
rect 205102 277618 240546 277854
rect 240782 277618 240866 277854
rect 241102 277618 276546 277854
rect 276782 277618 276866 277854
rect 277102 277618 312546 277854
rect 312782 277618 312866 277854
rect 313102 277618 348546 277854
rect 348782 277618 348866 277854
rect 349102 277618 384546 277854
rect 384782 277618 384866 277854
rect 385102 277618 420546 277854
rect 420782 277618 420866 277854
rect 421102 277618 456546 277854
rect 456782 277618 456866 277854
rect 457102 277618 492546 277854
rect 492782 277618 492866 277854
rect 493102 277618 528546 277854
rect 528782 277618 528866 277854
rect 529102 277618 564546 277854
rect 564782 277618 564866 277854
rect 565102 277618 591102 277854
rect 591338 277618 591422 277854
rect 591658 277618 592650 277854
rect -8726 277586 592650 277618
rect -8726 274454 592650 274486
rect -8726 274218 -6774 274454
rect -6538 274218 -6454 274454
rect -6218 274218 20826 274454
rect 21062 274218 21146 274454
rect 21382 274218 56826 274454
rect 57062 274218 57146 274454
rect 57382 274218 92826 274454
rect 93062 274218 93146 274454
rect 93382 274218 128826 274454
rect 129062 274218 129146 274454
rect 129382 274218 164826 274454
rect 165062 274218 165146 274454
rect 165382 274218 200826 274454
rect 201062 274218 201146 274454
rect 201382 274218 236826 274454
rect 237062 274218 237146 274454
rect 237382 274218 272826 274454
rect 273062 274218 273146 274454
rect 273382 274218 308826 274454
rect 309062 274218 309146 274454
rect 309382 274218 344826 274454
rect 345062 274218 345146 274454
rect 345382 274218 380826 274454
rect 381062 274218 381146 274454
rect 381382 274218 416826 274454
rect 417062 274218 417146 274454
rect 417382 274218 452826 274454
rect 453062 274218 453146 274454
rect 453382 274218 488826 274454
rect 489062 274218 489146 274454
rect 489382 274218 524826 274454
rect 525062 274218 525146 274454
rect 525382 274218 560826 274454
rect 561062 274218 561146 274454
rect 561382 274218 590142 274454
rect 590378 274218 590462 274454
rect 590698 274218 592650 274454
rect -8726 274134 592650 274218
rect -8726 273898 -6774 274134
rect -6538 273898 -6454 274134
rect -6218 273898 20826 274134
rect 21062 273898 21146 274134
rect 21382 273898 56826 274134
rect 57062 273898 57146 274134
rect 57382 273898 92826 274134
rect 93062 273898 93146 274134
rect 93382 273898 128826 274134
rect 129062 273898 129146 274134
rect 129382 273898 164826 274134
rect 165062 273898 165146 274134
rect 165382 273898 200826 274134
rect 201062 273898 201146 274134
rect 201382 273898 236826 274134
rect 237062 273898 237146 274134
rect 237382 273898 272826 274134
rect 273062 273898 273146 274134
rect 273382 273898 308826 274134
rect 309062 273898 309146 274134
rect 309382 273898 344826 274134
rect 345062 273898 345146 274134
rect 345382 273898 380826 274134
rect 381062 273898 381146 274134
rect 381382 273898 416826 274134
rect 417062 273898 417146 274134
rect 417382 273898 452826 274134
rect 453062 273898 453146 274134
rect 453382 273898 488826 274134
rect 489062 273898 489146 274134
rect 489382 273898 524826 274134
rect 525062 273898 525146 274134
rect 525382 273898 560826 274134
rect 561062 273898 561146 274134
rect 561382 273898 590142 274134
rect 590378 273898 590462 274134
rect 590698 273898 592650 274134
rect -8726 273866 592650 273898
rect -8726 270734 592650 270766
rect -8726 270498 -5814 270734
rect -5578 270498 -5494 270734
rect -5258 270498 17106 270734
rect 17342 270498 17426 270734
rect 17662 270498 53106 270734
rect 53342 270498 53426 270734
rect 53662 270498 89106 270734
rect 89342 270498 89426 270734
rect 89662 270498 125106 270734
rect 125342 270498 125426 270734
rect 125662 270498 161106 270734
rect 161342 270498 161426 270734
rect 161662 270498 197106 270734
rect 197342 270498 197426 270734
rect 197662 270498 233106 270734
rect 233342 270498 233426 270734
rect 233662 270498 269106 270734
rect 269342 270498 269426 270734
rect 269662 270498 305106 270734
rect 305342 270498 305426 270734
rect 305662 270498 341106 270734
rect 341342 270498 341426 270734
rect 341662 270498 377106 270734
rect 377342 270498 377426 270734
rect 377662 270498 413106 270734
rect 413342 270498 413426 270734
rect 413662 270498 449106 270734
rect 449342 270498 449426 270734
rect 449662 270498 485106 270734
rect 485342 270498 485426 270734
rect 485662 270498 521106 270734
rect 521342 270498 521426 270734
rect 521662 270498 557106 270734
rect 557342 270498 557426 270734
rect 557662 270498 589182 270734
rect 589418 270498 589502 270734
rect 589738 270498 592650 270734
rect -8726 270414 592650 270498
rect -8726 270178 -5814 270414
rect -5578 270178 -5494 270414
rect -5258 270178 17106 270414
rect 17342 270178 17426 270414
rect 17662 270178 53106 270414
rect 53342 270178 53426 270414
rect 53662 270178 89106 270414
rect 89342 270178 89426 270414
rect 89662 270178 125106 270414
rect 125342 270178 125426 270414
rect 125662 270178 161106 270414
rect 161342 270178 161426 270414
rect 161662 270178 197106 270414
rect 197342 270178 197426 270414
rect 197662 270178 233106 270414
rect 233342 270178 233426 270414
rect 233662 270178 269106 270414
rect 269342 270178 269426 270414
rect 269662 270178 305106 270414
rect 305342 270178 305426 270414
rect 305662 270178 341106 270414
rect 341342 270178 341426 270414
rect 341662 270178 377106 270414
rect 377342 270178 377426 270414
rect 377662 270178 413106 270414
rect 413342 270178 413426 270414
rect 413662 270178 449106 270414
rect 449342 270178 449426 270414
rect 449662 270178 485106 270414
rect 485342 270178 485426 270414
rect 485662 270178 521106 270414
rect 521342 270178 521426 270414
rect 521662 270178 557106 270414
rect 557342 270178 557426 270414
rect 557662 270178 589182 270414
rect 589418 270178 589502 270414
rect 589738 270178 592650 270414
rect -8726 270146 592650 270178
rect -8726 267014 592650 267046
rect -8726 266778 -4854 267014
rect -4618 266778 -4534 267014
rect -4298 266778 13386 267014
rect 13622 266778 13706 267014
rect 13942 266778 49386 267014
rect 49622 266778 49706 267014
rect 49942 266778 85386 267014
rect 85622 266778 85706 267014
rect 85942 266778 121386 267014
rect 121622 266778 121706 267014
rect 121942 266778 157386 267014
rect 157622 266778 157706 267014
rect 157942 266778 193386 267014
rect 193622 266778 193706 267014
rect 193942 266778 229386 267014
rect 229622 266778 229706 267014
rect 229942 266778 265386 267014
rect 265622 266778 265706 267014
rect 265942 266778 301386 267014
rect 301622 266778 301706 267014
rect 301942 266778 337386 267014
rect 337622 266778 337706 267014
rect 337942 266778 373386 267014
rect 373622 266778 373706 267014
rect 373942 266778 409386 267014
rect 409622 266778 409706 267014
rect 409942 266778 445386 267014
rect 445622 266778 445706 267014
rect 445942 266778 481386 267014
rect 481622 266778 481706 267014
rect 481942 266778 517386 267014
rect 517622 266778 517706 267014
rect 517942 266778 553386 267014
rect 553622 266778 553706 267014
rect 553942 266778 588222 267014
rect 588458 266778 588542 267014
rect 588778 266778 592650 267014
rect -8726 266694 592650 266778
rect -8726 266458 -4854 266694
rect -4618 266458 -4534 266694
rect -4298 266458 13386 266694
rect 13622 266458 13706 266694
rect 13942 266458 49386 266694
rect 49622 266458 49706 266694
rect 49942 266458 85386 266694
rect 85622 266458 85706 266694
rect 85942 266458 121386 266694
rect 121622 266458 121706 266694
rect 121942 266458 157386 266694
rect 157622 266458 157706 266694
rect 157942 266458 193386 266694
rect 193622 266458 193706 266694
rect 193942 266458 229386 266694
rect 229622 266458 229706 266694
rect 229942 266458 265386 266694
rect 265622 266458 265706 266694
rect 265942 266458 301386 266694
rect 301622 266458 301706 266694
rect 301942 266458 337386 266694
rect 337622 266458 337706 266694
rect 337942 266458 373386 266694
rect 373622 266458 373706 266694
rect 373942 266458 409386 266694
rect 409622 266458 409706 266694
rect 409942 266458 445386 266694
rect 445622 266458 445706 266694
rect 445942 266458 481386 266694
rect 481622 266458 481706 266694
rect 481942 266458 517386 266694
rect 517622 266458 517706 266694
rect 517942 266458 553386 266694
rect 553622 266458 553706 266694
rect 553942 266458 588222 266694
rect 588458 266458 588542 266694
rect 588778 266458 592650 266694
rect -8726 266426 592650 266458
rect -8726 263294 592650 263326
rect -8726 263058 -3894 263294
rect -3658 263058 -3574 263294
rect -3338 263058 9666 263294
rect 9902 263058 9986 263294
rect 10222 263058 45666 263294
rect 45902 263058 45986 263294
rect 46222 263058 81666 263294
rect 81902 263058 81986 263294
rect 82222 263058 117666 263294
rect 117902 263058 117986 263294
rect 118222 263058 153666 263294
rect 153902 263058 153986 263294
rect 154222 263058 189666 263294
rect 189902 263058 189986 263294
rect 190222 263058 225666 263294
rect 225902 263058 225986 263294
rect 226222 263058 261666 263294
rect 261902 263058 261986 263294
rect 262222 263058 297666 263294
rect 297902 263058 297986 263294
rect 298222 263058 333666 263294
rect 333902 263058 333986 263294
rect 334222 263058 369666 263294
rect 369902 263058 369986 263294
rect 370222 263058 405666 263294
rect 405902 263058 405986 263294
rect 406222 263058 441666 263294
rect 441902 263058 441986 263294
rect 442222 263058 477666 263294
rect 477902 263058 477986 263294
rect 478222 263058 513666 263294
rect 513902 263058 513986 263294
rect 514222 263058 549666 263294
rect 549902 263058 549986 263294
rect 550222 263058 587262 263294
rect 587498 263058 587582 263294
rect 587818 263058 592650 263294
rect -8726 262974 592650 263058
rect -8726 262738 -3894 262974
rect -3658 262738 -3574 262974
rect -3338 262738 9666 262974
rect 9902 262738 9986 262974
rect 10222 262738 45666 262974
rect 45902 262738 45986 262974
rect 46222 262738 81666 262974
rect 81902 262738 81986 262974
rect 82222 262738 117666 262974
rect 117902 262738 117986 262974
rect 118222 262738 153666 262974
rect 153902 262738 153986 262974
rect 154222 262738 189666 262974
rect 189902 262738 189986 262974
rect 190222 262738 225666 262974
rect 225902 262738 225986 262974
rect 226222 262738 261666 262974
rect 261902 262738 261986 262974
rect 262222 262738 297666 262974
rect 297902 262738 297986 262974
rect 298222 262738 333666 262974
rect 333902 262738 333986 262974
rect 334222 262738 369666 262974
rect 369902 262738 369986 262974
rect 370222 262738 405666 262974
rect 405902 262738 405986 262974
rect 406222 262738 441666 262974
rect 441902 262738 441986 262974
rect 442222 262738 477666 262974
rect 477902 262738 477986 262974
rect 478222 262738 513666 262974
rect 513902 262738 513986 262974
rect 514222 262738 549666 262974
rect 549902 262738 549986 262974
rect 550222 262738 587262 262974
rect 587498 262738 587582 262974
rect 587818 262738 592650 262974
rect -8726 262706 592650 262738
rect -8726 259574 592650 259606
rect -8726 259338 -2934 259574
rect -2698 259338 -2614 259574
rect -2378 259338 5946 259574
rect 6182 259338 6266 259574
rect 6502 259338 41946 259574
rect 42182 259338 42266 259574
rect 42502 259338 77946 259574
rect 78182 259338 78266 259574
rect 78502 259338 113946 259574
rect 114182 259338 114266 259574
rect 114502 259338 149946 259574
rect 150182 259338 150266 259574
rect 150502 259338 185946 259574
rect 186182 259338 186266 259574
rect 186502 259338 221946 259574
rect 222182 259338 222266 259574
rect 222502 259338 257946 259574
rect 258182 259338 258266 259574
rect 258502 259338 293946 259574
rect 294182 259338 294266 259574
rect 294502 259338 329946 259574
rect 330182 259338 330266 259574
rect 330502 259338 365946 259574
rect 366182 259338 366266 259574
rect 366502 259338 401946 259574
rect 402182 259338 402266 259574
rect 402502 259338 437946 259574
rect 438182 259338 438266 259574
rect 438502 259338 473946 259574
rect 474182 259338 474266 259574
rect 474502 259338 509946 259574
rect 510182 259338 510266 259574
rect 510502 259338 545946 259574
rect 546182 259338 546266 259574
rect 546502 259338 581946 259574
rect 582182 259338 582266 259574
rect 582502 259338 586302 259574
rect 586538 259338 586622 259574
rect 586858 259338 592650 259574
rect -8726 259254 592650 259338
rect -8726 259018 -2934 259254
rect -2698 259018 -2614 259254
rect -2378 259018 5946 259254
rect 6182 259018 6266 259254
rect 6502 259018 41946 259254
rect 42182 259018 42266 259254
rect 42502 259018 77946 259254
rect 78182 259018 78266 259254
rect 78502 259018 113946 259254
rect 114182 259018 114266 259254
rect 114502 259018 149946 259254
rect 150182 259018 150266 259254
rect 150502 259018 185946 259254
rect 186182 259018 186266 259254
rect 186502 259018 221946 259254
rect 222182 259018 222266 259254
rect 222502 259018 257946 259254
rect 258182 259018 258266 259254
rect 258502 259018 293946 259254
rect 294182 259018 294266 259254
rect 294502 259018 329946 259254
rect 330182 259018 330266 259254
rect 330502 259018 365946 259254
rect 366182 259018 366266 259254
rect 366502 259018 401946 259254
rect 402182 259018 402266 259254
rect 402502 259018 437946 259254
rect 438182 259018 438266 259254
rect 438502 259018 473946 259254
rect 474182 259018 474266 259254
rect 474502 259018 509946 259254
rect 510182 259018 510266 259254
rect 510502 259018 545946 259254
rect 546182 259018 546266 259254
rect 546502 259018 581946 259254
rect 582182 259018 582266 259254
rect 582502 259018 586302 259254
rect 586538 259018 586622 259254
rect 586858 259018 592650 259254
rect -8726 258986 592650 259018
rect -8726 255854 592650 255886
rect -8726 255618 -1974 255854
rect -1738 255618 -1654 255854
rect -1418 255618 2226 255854
rect 2462 255618 2546 255854
rect 2782 255618 38226 255854
rect 38462 255618 38546 255854
rect 38782 255618 74226 255854
rect 74462 255618 74546 255854
rect 74782 255618 110226 255854
rect 110462 255618 110546 255854
rect 110782 255618 146226 255854
rect 146462 255618 146546 255854
rect 146782 255618 182226 255854
rect 182462 255618 182546 255854
rect 182782 255618 218226 255854
rect 218462 255618 218546 255854
rect 218782 255618 254226 255854
rect 254462 255618 254546 255854
rect 254782 255618 290226 255854
rect 290462 255618 290546 255854
rect 290782 255618 326226 255854
rect 326462 255618 326546 255854
rect 326782 255618 362226 255854
rect 362462 255618 362546 255854
rect 362782 255618 398226 255854
rect 398462 255618 398546 255854
rect 398782 255618 434226 255854
rect 434462 255618 434546 255854
rect 434782 255618 470226 255854
rect 470462 255618 470546 255854
rect 470782 255618 506226 255854
rect 506462 255618 506546 255854
rect 506782 255618 542226 255854
rect 542462 255618 542546 255854
rect 542782 255618 578226 255854
rect 578462 255618 578546 255854
rect 578782 255618 585342 255854
rect 585578 255618 585662 255854
rect 585898 255618 592650 255854
rect -8726 255534 592650 255618
rect -8726 255298 -1974 255534
rect -1738 255298 -1654 255534
rect -1418 255298 2226 255534
rect 2462 255298 2546 255534
rect 2782 255298 38226 255534
rect 38462 255298 38546 255534
rect 38782 255298 74226 255534
rect 74462 255298 74546 255534
rect 74782 255298 110226 255534
rect 110462 255298 110546 255534
rect 110782 255298 146226 255534
rect 146462 255298 146546 255534
rect 146782 255298 182226 255534
rect 182462 255298 182546 255534
rect 182782 255298 218226 255534
rect 218462 255298 218546 255534
rect 218782 255298 254226 255534
rect 254462 255298 254546 255534
rect 254782 255298 290226 255534
rect 290462 255298 290546 255534
rect 290782 255298 326226 255534
rect 326462 255298 326546 255534
rect 326782 255298 362226 255534
rect 362462 255298 362546 255534
rect 362782 255298 398226 255534
rect 398462 255298 398546 255534
rect 398782 255298 434226 255534
rect 434462 255298 434546 255534
rect 434782 255298 470226 255534
rect 470462 255298 470546 255534
rect 470782 255298 506226 255534
rect 506462 255298 506546 255534
rect 506782 255298 542226 255534
rect 542462 255298 542546 255534
rect 542782 255298 578226 255534
rect 578462 255298 578546 255534
rect 578782 255298 585342 255534
rect 585578 255298 585662 255534
rect 585898 255298 592650 255534
rect -8726 255266 592650 255298
rect -8726 245894 592650 245926
rect -8726 245658 -8694 245894
rect -8458 245658 -8374 245894
rect -8138 245658 28266 245894
rect 28502 245658 28586 245894
rect 28822 245658 64266 245894
rect 64502 245658 64586 245894
rect 64822 245658 100266 245894
rect 100502 245658 100586 245894
rect 100822 245658 136266 245894
rect 136502 245658 136586 245894
rect 136822 245658 172266 245894
rect 172502 245658 172586 245894
rect 172822 245658 208266 245894
rect 208502 245658 208586 245894
rect 208822 245658 244266 245894
rect 244502 245658 244586 245894
rect 244822 245658 280266 245894
rect 280502 245658 280586 245894
rect 280822 245658 316266 245894
rect 316502 245658 316586 245894
rect 316822 245658 352266 245894
rect 352502 245658 352586 245894
rect 352822 245658 388266 245894
rect 388502 245658 388586 245894
rect 388822 245658 424266 245894
rect 424502 245658 424586 245894
rect 424822 245658 460266 245894
rect 460502 245658 460586 245894
rect 460822 245658 496266 245894
rect 496502 245658 496586 245894
rect 496822 245658 532266 245894
rect 532502 245658 532586 245894
rect 532822 245658 568266 245894
rect 568502 245658 568586 245894
rect 568822 245658 592062 245894
rect 592298 245658 592382 245894
rect 592618 245658 592650 245894
rect -8726 245574 592650 245658
rect -8726 245338 -8694 245574
rect -8458 245338 -8374 245574
rect -8138 245338 28266 245574
rect 28502 245338 28586 245574
rect 28822 245338 64266 245574
rect 64502 245338 64586 245574
rect 64822 245338 100266 245574
rect 100502 245338 100586 245574
rect 100822 245338 136266 245574
rect 136502 245338 136586 245574
rect 136822 245338 172266 245574
rect 172502 245338 172586 245574
rect 172822 245338 208266 245574
rect 208502 245338 208586 245574
rect 208822 245338 244266 245574
rect 244502 245338 244586 245574
rect 244822 245338 280266 245574
rect 280502 245338 280586 245574
rect 280822 245338 316266 245574
rect 316502 245338 316586 245574
rect 316822 245338 352266 245574
rect 352502 245338 352586 245574
rect 352822 245338 388266 245574
rect 388502 245338 388586 245574
rect 388822 245338 424266 245574
rect 424502 245338 424586 245574
rect 424822 245338 460266 245574
rect 460502 245338 460586 245574
rect 460822 245338 496266 245574
rect 496502 245338 496586 245574
rect 496822 245338 532266 245574
rect 532502 245338 532586 245574
rect 532822 245338 568266 245574
rect 568502 245338 568586 245574
rect 568822 245338 592062 245574
rect 592298 245338 592382 245574
rect 592618 245338 592650 245574
rect -8726 245306 592650 245338
rect -8726 242174 592650 242206
rect -8726 241938 -7734 242174
rect -7498 241938 -7414 242174
rect -7178 241938 24546 242174
rect 24782 241938 24866 242174
rect 25102 241938 60546 242174
rect 60782 241938 60866 242174
rect 61102 241938 96546 242174
rect 96782 241938 96866 242174
rect 97102 241938 132546 242174
rect 132782 241938 132866 242174
rect 133102 241938 168546 242174
rect 168782 241938 168866 242174
rect 169102 241938 204546 242174
rect 204782 241938 204866 242174
rect 205102 241938 240546 242174
rect 240782 241938 240866 242174
rect 241102 241938 276546 242174
rect 276782 241938 276866 242174
rect 277102 241938 312546 242174
rect 312782 241938 312866 242174
rect 313102 241938 348546 242174
rect 348782 241938 348866 242174
rect 349102 241938 384546 242174
rect 384782 241938 384866 242174
rect 385102 241938 420546 242174
rect 420782 241938 420866 242174
rect 421102 241938 456546 242174
rect 456782 241938 456866 242174
rect 457102 241938 492546 242174
rect 492782 241938 492866 242174
rect 493102 241938 528546 242174
rect 528782 241938 528866 242174
rect 529102 241938 564546 242174
rect 564782 241938 564866 242174
rect 565102 241938 591102 242174
rect 591338 241938 591422 242174
rect 591658 241938 592650 242174
rect -8726 241854 592650 241938
rect -8726 241618 -7734 241854
rect -7498 241618 -7414 241854
rect -7178 241618 24546 241854
rect 24782 241618 24866 241854
rect 25102 241618 60546 241854
rect 60782 241618 60866 241854
rect 61102 241618 96546 241854
rect 96782 241618 96866 241854
rect 97102 241618 132546 241854
rect 132782 241618 132866 241854
rect 133102 241618 168546 241854
rect 168782 241618 168866 241854
rect 169102 241618 204546 241854
rect 204782 241618 204866 241854
rect 205102 241618 240546 241854
rect 240782 241618 240866 241854
rect 241102 241618 276546 241854
rect 276782 241618 276866 241854
rect 277102 241618 312546 241854
rect 312782 241618 312866 241854
rect 313102 241618 348546 241854
rect 348782 241618 348866 241854
rect 349102 241618 384546 241854
rect 384782 241618 384866 241854
rect 385102 241618 420546 241854
rect 420782 241618 420866 241854
rect 421102 241618 456546 241854
rect 456782 241618 456866 241854
rect 457102 241618 492546 241854
rect 492782 241618 492866 241854
rect 493102 241618 528546 241854
rect 528782 241618 528866 241854
rect 529102 241618 564546 241854
rect 564782 241618 564866 241854
rect 565102 241618 591102 241854
rect 591338 241618 591422 241854
rect 591658 241618 592650 241854
rect -8726 241586 592650 241618
rect -8726 238454 592650 238486
rect -8726 238218 -6774 238454
rect -6538 238218 -6454 238454
rect -6218 238218 20826 238454
rect 21062 238218 21146 238454
rect 21382 238218 56826 238454
rect 57062 238218 57146 238454
rect 57382 238218 92826 238454
rect 93062 238218 93146 238454
rect 93382 238218 128826 238454
rect 129062 238218 129146 238454
rect 129382 238218 164826 238454
rect 165062 238218 165146 238454
rect 165382 238218 200826 238454
rect 201062 238218 201146 238454
rect 201382 238218 236826 238454
rect 237062 238218 237146 238454
rect 237382 238218 272826 238454
rect 273062 238218 273146 238454
rect 273382 238218 308826 238454
rect 309062 238218 309146 238454
rect 309382 238218 344826 238454
rect 345062 238218 345146 238454
rect 345382 238218 380826 238454
rect 381062 238218 381146 238454
rect 381382 238218 416826 238454
rect 417062 238218 417146 238454
rect 417382 238218 452826 238454
rect 453062 238218 453146 238454
rect 453382 238218 488826 238454
rect 489062 238218 489146 238454
rect 489382 238218 524826 238454
rect 525062 238218 525146 238454
rect 525382 238218 560826 238454
rect 561062 238218 561146 238454
rect 561382 238218 590142 238454
rect 590378 238218 590462 238454
rect 590698 238218 592650 238454
rect -8726 238134 592650 238218
rect -8726 237898 -6774 238134
rect -6538 237898 -6454 238134
rect -6218 237898 20826 238134
rect 21062 237898 21146 238134
rect 21382 237898 56826 238134
rect 57062 237898 57146 238134
rect 57382 237898 92826 238134
rect 93062 237898 93146 238134
rect 93382 237898 128826 238134
rect 129062 237898 129146 238134
rect 129382 237898 164826 238134
rect 165062 237898 165146 238134
rect 165382 237898 200826 238134
rect 201062 237898 201146 238134
rect 201382 237898 236826 238134
rect 237062 237898 237146 238134
rect 237382 237898 272826 238134
rect 273062 237898 273146 238134
rect 273382 237898 308826 238134
rect 309062 237898 309146 238134
rect 309382 237898 344826 238134
rect 345062 237898 345146 238134
rect 345382 237898 380826 238134
rect 381062 237898 381146 238134
rect 381382 237898 416826 238134
rect 417062 237898 417146 238134
rect 417382 237898 452826 238134
rect 453062 237898 453146 238134
rect 453382 237898 488826 238134
rect 489062 237898 489146 238134
rect 489382 237898 524826 238134
rect 525062 237898 525146 238134
rect 525382 237898 560826 238134
rect 561062 237898 561146 238134
rect 561382 237898 590142 238134
rect 590378 237898 590462 238134
rect 590698 237898 592650 238134
rect -8726 237866 592650 237898
rect -8726 234734 592650 234766
rect -8726 234498 -5814 234734
rect -5578 234498 -5494 234734
rect -5258 234498 17106 234734
rect 17342 234498 17426 234734
rect 17662 234498 53106 234734
rect 53342 234498 53426 234734
rect 53662 234498 89106 234734
rect 89342 234498 89426 234734
rect 89662 234498 125106 234734
rect 125342 234498 125426 234734
rect 125662 234498 161106 234734
rect 161342 234498 161426 234734
rect 161662 234498 197106 234734
rect 197342 234498 197426 234734
rect 197662 234498 233106 234734
rect 233342 234498 233426 234734
rect 233662 234498 269106 234734
rect 269342 234498 269426 234734
rect 269662 234498 305106 234734
rect 305342 234498 305426 234734
rect 305662 234498 341106 234734
rect 341342 234498 341426 234734
rect 341662 234498 377106 234734
rect 377342 234498 377426 234734
rect 377662 234498 413106 234734
rect 413342 234498 413426 234734
rect 413662 234498 449106 234734
rect 449342 234498 449426 234734
rect 449662 234498 485106 234734
rect 485342 234498 485426 234734
rect 485662 234498 521106 234734
rect 521342 234498 521426 234734
rect 521662 234498 557106 234734
rect 557342 234498 557426 234734
rect 557662 234498 589182 234734
rect 589418 234498 589502 234734
rect 589738 234498 592650 234734
rect -8726 234414 592650 234498
rect -8726 234178 -5814 234414
rect -5578 234178 -5494 234414
rect -5258 234178 17106 234414
rect 17342 234178 17426 234414
rect 17662 234178 53106 234414
rect 53342 234178 53426 234414
rect 53662 234178 89106 234414
rect 89342 234178 89426 234414
rect 89662 234178 125106 234414
rect 125342 234178 125426 234414
rect 125662 234178 161106 234414
rect 161342 234178 161426 234414
rect 161662 234178 197106 234414
rect 197342 234178 197426 234414
rect 197662 234178 233106 234414
rect 233342 234178 233426 234414
rect 233662 234178 269106 234414
rect 269342 234178 269426 234414
rect 269662 234178 305106 234414
rect 305342 234178 305426 234414
rect 305662 234178 341106 234414
rect 341342 234178 341426 234414
rect 341662 234178 377106 234414
rect 377342 234178 377426 234414
rect 377662 234178 413106 234414
rect 413342 234178 413426 234414
rect 413662 234178 449106 234414
rect 449342 234178 449426 234414
rect 449662 234178 485106 234414
rect 485342 234178 485426 234414
rect 485662 234178 521106 234414
rect 521342 234178 521426 234414
rect 521662 234178 557106 234414
rect 557342 234178 557426 234414
rect 557662 234178 589182 234414
rect 589418 234178 589502 234414
rect 589738 234178 592650 234414
rect -8726 234146 592650 234178
rect -8726 231014 592650 231046
rect -8726 230778 -4854 231014
rect -4618 230778 -4534 231014
rect -4298 230778 13386 231014
rect 13622 230778 13706 231014
rect 13942 230778 49386 231014
rect 49622 230778 49706 231014
rect 49942 230778 85386 231014
rect 85622 230778 85706 231014
rect 85942 230778 121386 231014
rect 121622 230778 121706 231014
rect 121942 230778 157386 231014
rect 157622 230778 157706 231014
rect 157942 230778 193386 231014
rect 193622 230778 193706 231014
rect 193942 230778 229386 231014
rect 229622 230778 229706 231014
rect 229942 230778 265386 231014
rect 265622 230778 265706 231014
rect 265942 230778 301386 231014
rect 301622 230778 301706 231014
rect 301942 230778 337386 231014
rect 337622 230778 337706 231014
rect 337942 230778 373386 231014
rect 373622 230778 373706 231014
rect 373942 230778 409386 231014
rect 409622 230778 409706 231014
rect 409942 230778 445386 231014
rect 445622 230778 445706 231014
rect 445942 230778 481386 231014
rect 481622 230778 481706 231014
rect 481942 230778 517386 231014
rect 517622 230778 517706 231014
rect 517942 230778 553386 231014
rect 553622 230778 553706 231014
rect 553942 230778 588222 231014
rect 588458 230778 588542 231014
rect 588778 230778 592650 231014
rect -8726 230694 592650 230778
rect -8726 230458 -4854 230694
rect -4618 230458 -4534 230694
rect -4298 230458 13386 230694
rect 13622 230458 13706 230694
rect 13942 230458 49386 230694
rect 49622 230458 49706 230694
rect 49942 230458 85386 230694
rect 85622 230458 85706 230694
rect 85942 230458 121386 230694
rect 121622 230458 121706 230694
rect 121942 230458 157386 230694
rect 157622 230458 157706 230694
rect 157942 230458 193386 230694
rect 193622 230458 193706 230694
rect 193942 230458 229386 230694
rect 229622 230458 229706 230694
rect 229942 230458 265386 230694
rect 265622 230458 265706 230694
rect 265942 230458 301386 230694
rect 301622 230458 301706 230694
rect 301942 230458 337386 230694
rect 337622 230458 337706 230694
rect 337942 230458 373386 230694
rect 373622 230458 373706 230694
rect 373942 230458 409386 230694
rect 409622 230458 409706 230694
rect 409942 230458 445386 230694
rect 445622 230458 445706 230694
rect 445942 230458 481386 230694
rect 481622 230458 481706 230694
rect 481942 230458 517386 230694
rect 517622 230458 517706 230694
rect 517942 230458 553386 230694
rect 553622 230458 553706 230694
rect 553942 230458 588222 230694
rect 588458 230458 588542 230694
rect 588778 230458 592650 230694
rect -8726 230426 592650 230458
rect -8726 227294 592650 227326
rect -8726 227058 -3894 227294
rect -3658 227058 -3574 227294
rect -3338 227058 9666 227294
rect 9902 227058 9986 227294
rect 10222 227058 45666 227294
rect 45902 227058 45986 227294
rect 46222 227058 81666 227294
rect 81902 227058 81986 227294
rect 82222 227058 117666 227294
rect 117902 227058 117986 227294
rect 118222 227058 153666 227294
rect 153902 227058 153986 227294
rect 154222 227058 189666 227294
rect 189902 227058 189986 227294
rect 190222 227058 225666 227294
rect 225902 227058 225986 227294
rect 226222 227058 261666 227294
rect 261902 227058 261986 227294
rect 262222 227058 297666 227294
rect 297902 227058 297986 227294
rect 298222 227058 333666 227294
rect 333902 227058 333986 227294
rect 334222 227058 369666 227294
rect 369902 227058 369986 227294
rect 370222 227058 405666 227294
rect 405902 227058 405986 227294
rect 406222 227058 441666 227294
rect 441902 227058 441986 227294
rect 442222 227058 477666 227294
rect 477902 227058 477986 227294
rect 478222 227058 513666 227294
rect 513902 227058 513986 227294
rect 514222 227058 549666 227294
rect 549902 227058 549986 227294
rect 550222 227058 587262 227294
rect 587498 227058 587582 227294
rect 587818 227058 592650 227294
rect -8726 226974 592650 227058
rect -8726 226738 -3894 226974
rect -3658 226738 -3574 226974
rect -3338 226738 9666 226974
rect 9902 226738 9986 226974
rect 10222 226738 45666 226974
rect 45902 226738 45986 226974
rect 46222 226738 81666 226974
rect 81902 226738 81986 226974
rect 82222 226738 117666 226974
rect 117902 226738 117986 226974
rect 118222 226738 153666 226974
rect 153902 226738 153986 226974
rect 154222 226738 189666 226974
rect 189902 226738 189986 226974
rect 190222 226738 225666 226974
rect 225902 226738 225986 226974
rect 226222 226738 261666 226974
rect 261902 226738 261986 226974
rect 262222 226738 297666 226974
rect 297902 226738 297986 226974
rect 298222 226738 333666 226974
rect 333902 226738 333986 226974
rect 334222 226738 369666 226974
rect 369902 226738 369986 226974
rect 370222 226738 405666 226974
rect 405902 226738 405986 226974
rect 406222 226738 441666 226974
rect 441902 226738 441986 226974
rect 442222 226738 477666 226974
rect 477902 226738 477986 226974
rect 478222 226738 513666 226974
rect 513902 226738 513986 226974
rect 514222 226738 549666 226974
rect 549902 226738 549986 226974
rect 550222 226738 587262 226974
rect 587498 226738 587582 226974
rect 587818 226738 592650 226974
rect -8726 226706 592650 226738
rect -8726 223574 592650 223606
rect -8726 223338 -2934 223574
rect -2698 223338 -2614 223574
rect -2378 223338 5946 223574
rect 6182 223338 6266 223574
rect 6502 223338 41946 223574
rect 42182 223338 42266 223574
rect 42502 223338 77946 223574
rect 78182 223338 78266 223574
rect 78502 223338 113946 223574
rect 114182 223338 114266 223574
rect 114502 223338 149946 223574
rect 150182 223338 150266 223574
rect 150502 223338 185946 223574
rect 186182 223338 186266 223574
rect 186502 223338 221946 223574
rect 222182 223338 222266 223574
rect 222502 223338 257946 223574
rect 258182 223338 258266 223574
rect 258502 223338 293946 223574
rect 294182 223338 294266 223574
rect 294502 223338 329946 223574
rect 330182 223338 330266 223574
rect 330502 223338 365946 223574
rect 366182 223338 366266 223574
rect 366502 223338 401946 223574
rect 402182 223338 402266 223574
rect 402502 223338 437946 223574
rect 438182 223338 438266 223574
rect 438502 223338 473946 223574
rect 474182 223338 474266 223574
rect 474502 223338 509946 223574
rect 510182 223338 510266 223574
rect 510502 223338 545946 223574
rect 546182 223338 546266 223574
rect 546502 223338 581946 223574
rect 582182 223338 582266 223574
rect 582502 223338 586302 223574
rect 586538 223338 586622 223574
rect 586858 223338 592650 223574
rect -8726 223254 592650 223338
rect -8726 223018 -2934 223254
rect -2698 223018 -2614 223254
rect -2378 223018 5946 223254
rect 6182 223018 6266 223254
rect 6502 223018 41946 223254
rect 42182 223018 42266 223254
rect 42502 223018 77946 223254
rect 78182 223018 78266 223254
rect 78502 223018 113946 223254
rect 114182 223018 114266 223254
rect 114502 223018 149946 223254
rect 150182 223018 150266 223254
rect 150502 223018 185946 223254
rect 186182 223018 186266 223254
rect 186502 223018 221946 223254
rect 222182 223018 222266 223254
rect 222502 223018 257946 223254
rect 258182 223018 258266 223254
rect 258502 223018 293946 223254
rect 294182 223018 294266 223254
rect 294502 223018 329946 223254
rect 330182 223018 330266 223254
rect 330502 223018 365946 223254
rect 366182 223018 366266 223254
rect 366502 223018 401946 223254
rect 402182 223018 402266 223254
rect 402502 223018 437946 223254
rect 438182 223018 438266 223254
rect 438502 223018 473946 223254
rect 474182 223018 474266 223254
rect 474502 223018 509946 223254
rect 510182 223018 510266 223254
rect 510502 223018 545946 223254
rect 546182 223018 546266 223254
rect 546502 223018 581946 223254
rect 582182 223018 582266 223254
rect 582502 223018 586302 223254
rect 586538 223018 586622 223254
rect 586858 223018 592650 223254
rect -8726 222986 592650 223018
rect -8726 219854 592650 219886
rect -8726 219618 -1974 219854
rect -1738 219618 -1654 219854
rect -1418 219618 2226 219854
rect 2462 219618 2546 219854
rect 2782 219618 38226 219854
rect 38462 219618 38546 219854
rect 38782 219618 74226 219854
rect 74462 219618 74546 219854
rect 74782 219618 110226 219854
rect 110462 219618 110546 219854
rect 110782 219618 146226 219854
rect 146462 219618 146546 219854
rect 146782 219618 182226 219854
rect 182462 219618 182546 219854
rect 182782 219618 218226 219854
rect 218462 219618 218546 219854
rect 218782 219618 254226 219854
rect 254462 219618 254546 219854
rect 254782 219618 290226 219854
rect 290462 219618 290546 219854
rect 290782 219618 326226 219854
rect 326462 219618 326546 219854
rect 326782 219618 362226 219854
rect 362462 219618 362546 219854
rect 362782 219618 398226 219854
rect 398462 219618 398546 219854
rect 398782 219618 434226 219854
rect 434462 219618 434546 219854
rect 434782 219618 470226 219854
rect 470462 219618 470546 219854
rect 470782 219618 506226 219854
rect 506462 219618 506546 219854
rect 506782 219618 542226 219854
rect 542462 219618 542546 219854
rect 542782 219618 578226 219854
rect 578462 219618 578546 219854
rect 578782 219618 585342 219854
rect 585578 219618 585662 219854
rect 585898 219618 592650 219854
rect -8726 219534 592650 219618
rect -8726 219298 -1974 219534
rect -1738 219298 -1654 219534
rect -1418 219298 2226 219534
rect 2462 219298 2546 219534
rect 2782 219298 38226 219534
rect 38462 219298 38546 219534
rect 38782 219298 74226 219534
rect 74462 219298 74546 219534
rect 74782 219298 110226 219534
rect 110462 219298 110546 219534
rect 110782 219298 146226 219534
rect 146462 219298 146546 219534
rect 146782 219298 182226 219534
rect 182462 219298 182546 219534
rect 182782 219298 218226 219534
rect 218462 219298 218546 219534
rect 218782 219298 254226 219534
rect 254462 219298 254546 219534
rect 254782 219298 290226 219534
rect 290462 219298 290546 219534
rect 290782 219298 326226 219534
rect 326462 219298 326546 219534
rect 326782 219298 362226 219534
rect 362462 219298 362546 219534
rect 362782 219298 398226 219534
rect 398462 219298 398546 219534
rect 398782 219298 434226 219534
rect 434462 219298 434546 219534
rect 434782 219298 470226 219534
rect 470462 219298 470546 219534
rect 470782 219298 506226 219534
rect 506462 219298 506546 219534
rect 506782 219298 542226 219534
rect 542462 219298 542546 219534
rect 542782 219298 578226 219534
rect 578462 219298 578546 219534
rect 578782 219298 585342 219534
rect 585578 219298 585662 219534
rect 585898 219298 592650 219534
rect -8726 219266 592650 219298
rect -8726 209894 592650 209926
rect -8726 209658 -8694 209894
rect -8458 209658 -8374 209894
rect -8138 209658 28266 209894
rect 28502 209658 28586 209894
rect 28822 209658 64266 209894
rect 64502 209658 64586 209894
rect 64822 209658 100266 209894
rect 100502 209658 100586 209894
rect 100822 209658 136266 209894
rect 136502 209658 136586 209894
rect 136822 209658 172266 209894
rect 172502 209658 172586 209894
rect 172822 209658 208266 209894
rect 208502 209658 208586 209894
rect 208822 209658 244266 209894
rect 244502 209658 244586 209894
rect 244822 209658 280266 209894
rect 280502 209658 280586 209894
rect 280822 209658 316266 209894
rect 316502 209658 316586 209894
rect 316822 209658 352266 209894
rect 352502 209658 352586 209894
rect 352822 209658 388266 209894
rect 388502 209658 388586 209894
rect 388822 209658 424266 209894
rect 424502 209658 424586 209894
rect 424822 209658 460266 209894
rect 460502 209658 460586 209894
rect 460822 209658 496266 209894
rect 496502 209658 496586 209894
rect 496822 209658 532266 209894
rect 532502 209658 532586 209894
rect 532822 209658 568266 209894
rect 568502 209658 568586 209894
rect 568822 209658 592062 209894
rect 592298 209658 592382 209894
rect 592618 209658 592650 209894
rect -8726 209574 592650 209658
rect -8726 209338 -8694 209574
rect -8458 209338 -8374 209574
rect -8138 209338 28266 209574
rect 28502 209338 28586 209574
rect 28822 209338 64266 209574
rect 64502 209338 64586 209574
rect 64822 209338 100266 209574
rect 100502 209338 100586 209574
rect 100822 209338 136266 209574
rect 136502 209338 136586 209574
rect 136822 209338 172266 209574
rect 172502 209338 172586 209574
rect 172822 209338 208266 209574
rect 208502 209338 208586 209574
rect 208822 209338 244266 209574
rect 244502 209338 244586 209574
rect 244822 209338 280266 209574
rect 280502 209338 280586 209574
rect 280822 209338 316266 209574
rect 316502 209338 316586 209574
rect 316822 209338 352266 209574
rect 352502 209338 352586 209574
rect 352822 209338 388266 209574
rect 388502 209338 388586 209574
rect 388822 209338 424266 209574
rect 424502 209338 424586 209574
rect 424822 209338 460266 209574
rect 460502 209338 460586 209574
rect 460822 209338 496266 209574
rect 496502 209338 496586 209574
rect 496822 209338 532266 209574
rect 532502 209338 532586 209574
rect 532822 209338 568266 209574
rect 568502 209338 568586 209574
rect 568822 209338 592062 209574
rect 592298 209338 592382 209574
rect 592618 209338 592650 209574
rect -8726 209306 592650 209338
rect -8726 206174 592650 206206
rect -8726 205938 -7734 206174
rect -7498 205938 -7414 206174
rect -7178 205938 24546 206174
rect 24782 205938 24866 206174
rect 25102 205938 60546 206174
rect 60782 205938 60866 206174
rect 61102 205938 96546 206174
rect 96782 205938 96866 206174
rect 97102 205938 132546 206174
rect 132782 205938 132866 206174
rect 133102 205938 168546 206174
rect 168782 205938 168866 206174
rect 169102 205938 204546 206174
rect 204782 205938 204866 206174
rect 205102 205938 240546 206174
rect 240782 205938 240866 206174
rect 241102 205938 276546 206174
rect 276782 205938 276866 206174
rect 277102 205938 312546 206174
rect 312782 205938 312866 206174
rect 313102 205938 348546 206174
rect 348782 205938 348866 206174
rect 349102 205938 384546 206174
rect 384782 205938 384866 206174
rect 385102 205938 420546 206174
rect 420782 205938 420866 206174
rect 421102 205938 456546 206174
rect 456782 205938 456866 206174
rect 457102 205938 492546 206174
rect 492782 205938 492866 206174
rect 493102 205938 528546 206174
rect 528782 205938 528866 206174
rect 529102 205938 564546 206174
rect 564782 205938 564866 206174
rect 565102 205938 591102 206174
rect 591338 205938 591422 206174
rect 591658 205938 592650 206174
rect -8726 205854 592650 205938
rect -8726 205618 -7734 205854
rect -7498 205618 -7414 205854
rect -7178 205618 24546 205854
rect 24782 205618 24866 205854
rect 25102 205618 60546 205854
rect 60782 205618 60866 205854
rect 61102 205618 96546 205854
rect 96782 205618 96866 205854
rect 97102 205618 132546 205854
rect 132782 205618 132866 205854
rect 133102 205618 168546 205854
rect 168782 205618 168866 205854
rect 169102 205618 204546 205854
rect 204782 205618 204866 205854
rect 205102 205618 240546 205854
rect 240782 205618 240866 205854
rect 241102 205618 276546 205854
rect 276782 205618 276866 205854
rect 277102 205618 312546 205854
rect 312782 205618 312866 205854
rect 313102 205618 348546 205854
rect 348782 205618 348866 205854
rect 349102 205618 384546 205854
rect 384782 205618 384866 205854
rect 385102 205618 420546 205854
rect 420782 205618 420866 205854
rect 421102 205618 456546 205854
rect 456782 205618 456866 205854
rect 457102 205618 492546 205854
rect 492782 205618 492866 205854
rect 493102 205618 528546 205854
rect 528782 205618 528866 205854
rect 529102 205618 564546 205854
rect 564782 205618 564866 205854
rect 565102 205618 591102 205854
rect 591338 205618 591422 205854
rect 591658 205618 592650 205854
rect -8726 205586 592650 205618
rect -8726 202454 592650 202486
rect -8726 202218 -6774 202454
rect -6538 202218 -6454 202454
rect -6218 202218 20826 202454
rect 21062 202218 21146 202454
rect 21382 202218 56826 202454
rect 57062 202218 57146 202454
rect 57382 202218 92826 202454
rect 93062 202218 93146 202454
rect 93382 202218 128826 202454
rect 129062 202218 129146 202454
rect 129382 202218 164826 202454
rect 165062 202218 165146 202454
rect 165382 202218 200826 202454
rect 201062 202218 201146 202454
rect 201382 202218 236826 202454
rect 237062 202218 237146 202454
rect 237382 202218 272826 202454
rect 273062 202218 273146 202454
rect 273382 202218 308826 202454
rect 309062 202218 309146 202454
rect 309382 202218 344826 202454
rect 345062 202218 345146 202454
rect 345382 202218 380826 202454
rect 381062 202218 381146 202454
rect 381382 202218 416826 202454
rect 417062 202218 417146 202454
rect 417382 202218 452826 202454
rect 453062 202218 453146 202454
rect 453382 202218 488826 202454
rect 489062 202218 489146 202454
rect 489382 202218 524826 202454
rect 525062 202218 525146 202454
rect 525382 202218 560826 202454
rect 561062 202218 561146 202454
rect 561382 202218 590142 202454
rect 590378 202218 590462 202454
rect 590698 202218 592650 202454
rect -8726 202134 592650 202218
rect -8726 201898 -6774 202134
rect -6538 201898 -6454 202134
rect -6218 201898 20826 202134
rect 21062 201898 21146 202134
rect 21382 201898 56826 202134
rect 57062 201898 57146 202134
rect 57382 201898 92826 202134
rect 93062 201898 93146 202134
rect 93382 201898 128826 202134
rect 129062 201898 129146 202134
rect 129382 201898 164826 202134
rect 165062 201898 165146 202134
rect 165382 201898 200826 202134
rect 201062 201898 201146 202134
rect 201382 201898 236826 202134
rect 237062 201898 237146 202134
rect 237382 201898 272826 202134
rect 273062 201898 273146 202134
rect 273382 201898 308826 202134
rect 309062 201898 309146 202134
rect 309382 201898 344826 202134
rect 345062 201898 345146 202134
rect 345382 201898 380826 202134
rect 381062 201898 381146 202134
rect 381382 201898 416826 202134
rect 417062 201898 417146 202134
rect 417382 201898 452826 202134
rect 453062 201898 453146 202134
rect 453382 201898 488826 202134
rect 489062 201898 489146 202134
rect 489382 201898 524826 202134
rect 525062 201898 525146 202134
rect 525382 201898 560826 202134
rect 561062 201898 561146 202134
rect 561382 201898 590142 202134
rect 590378 201898 590462 202134
rect 590698 201898 592650 202134
rect -8726 201866 592650 201898
rect -8726 198734 592650 198766
rect -8726 198498 -5814 198734
rect -5578 198498 -5494 198734
rect -5258 198498 17106 198734
rect 17342 198498 17426 198734
rect 17662 198498 53106 198734
rect 53342 198498 53426 198734
rect 53662 198498 89106 198734
rect 89342 198498 89426 198734
rect 89662 198498 125106 198734
rect 125342 198498 125426 198734
rect 125662 198498 161106 198734
rect 161342 198498 161426 198734
rect 161662 198498 197106 198734
rect 197342 198498 197426 198734
rect 197662 198498 233106 198734
rect 233342 198498 233426 198734
rect 233662 198498 269106 198734
rect 269342 198498 269426 198734
rect 269662 198498 305106 198734
rect 305342 198498 305426 198734
rect 305662 198498 341106 198734
rect 341342 198498 341426 198734
rect 341662 198498 377106 198734
rect 377342 198498 377426 198734
rect 377662 198498 413106 198734
rect 413342 198498 413426 198734
rect 413662 198498 449106 198734
rect 449342 198498 449426 198734
rect 449662 198498 485106 198734
rect 485342 198498 485426 198734
rect 485662 198498 521106 198734
rect 521342 198498 521426 198734
rect 521662 198498 557106 198734
rect 557342 198498 557426 198734
rect 557662 198498 589182 198734
rect 589418 198498 589502 198734
rect 589738 198498 592650 198734
rect -8726 198414 592650 198498
rect -8726 198178 -5814 198414
rect -5578 198178 -5494 198414
rect -5258 198178 17106 198414
rect 17342 198178 17426 198414
rect 17662 198178 53106 198414
rect 53342 198178 53426 198414
rect 53662 198178 89106 198414
rect 89342 198178 89426 198414
rect 89662 198178 125106 198414
rect 125342 198178 125426 198414
rect 125662 198178 161106 198414
rect 161342 198178 161426 198414
rect 161662 198178 197106 198414
rect 197342 198178 197426 198414
rect 197662 198178 233106 198414
rect 233342 198178 233426 198414
rect 233662 198178 269106 198414
rect 269342 198178 269426 198414
rect 269662 198178 305106 198414
rect 305342 198178 305426 198414
rect 305662 198178 341106 198414
rect 341342 198178 341426 198414
rect 341662 198178 377106 198414
rect 377342 198178 377426 198414
rect 377662 198178 413106 198414
rect 413342 198178 413426 198414
rect 413662 198178 449106 198414
rect 449342 198178 449426 198414
rect 449662 198178 485106 198414
rect 485342 198178 485426 198414
rect 485662 198178 521106 198414
rect 521342 198178 521426 198414
rect 521662 198178 557106 198414
rect 557342 198178 557426 198414
rect 557662 198178 589182 198414
rect 589418 198178 589502 198414
rect 589738 198178 592650 198414
rect -8726 198146 592650 198178
rect -8726 195014 592650 195046
rect -8726 194778 -4854 195014
rect -4618 194778 -4534 195014
rect -4298 194778 13386 195014
rect 13622 194778 13706 195014
rect 13942 194778 49386 195014
rect 49622 194778 49706 195014
rect 49942 194778 85386 195014
rect 85622 194778 85706 195014
rect 85942 194778 121386 195014
rect 121622 194778 121706 195014
rect 121942 194778 157386 195014
rect 157622 194778 157706 195014
rect 157942 194778 193386 195014
rect 193622 194778 193706 195014
rect 193942 194778 229386 195014
rect 229622 194778 229706 195014
rect 229942 194778 265386 195014
rect 265622 194778 265706 195014
rect 265942 194778 301386 195014
rect 301622 194778 301706 195014
rect 301942 194778 337386 195014
rect 337622 194778 337706 195014
rect 337942 194778 373386 195014
rect 373622 194778 373706 195014
rect 373942 194778 409386 195014
rect 409622 194778 409706 195014
rect 409942 194778 445386 195014
rect 445622 194778 445706 195014
rect 445942 194778 481386 195014
rect 481622 194778 481706 195014
rect 481942 194778 517386 195014
rect 517622 194778 517706 195014
rect 517942 194778 553386 195014
rect 553622 194778 553706 195014
rect 553942 194778 588222 195014
rect 588458 194778 588542 195014
rect 588778 194778 592650 195014
rect -8726 194694 592650 194778
rect -8726 194458 -4854 194694
rect -4618 194458 -4534 194694
rect -4298 194458 13386 194694
rect 13622 194458 13706 194694
rect 13942 194458 49386 194694
rect 49622 194458 49706 194694
rect 49942 194458 85386 194694
rect 85622 194458 85706 194694
rect 85942 194458 121386 194694
rect 121622 194458 121706 194694
rect 121942 194458 157386 194694
rect 157622 194458 157706 194694
rect 157942 194458 193386 194694
rect 193622 194458 193706 194694
rect 193942 194458 229386 194694
rect 229622 194458 229706 194694
rect 229942 194458 265386 194694
rect 265622 194458 265706 194694
rect 265942 194458 301386 194694
rect 301622 194458 301706 194694
rect 301942 194458 337386 194694
rect 337622 194458 337706 194694
rect 337942 194458 373386 194694
rect 373622 194458 373706 194694
rect 373942 194458 409386 194694
rect 409622 194458 409706 194694
rect 409942 194458 445386 194694
rect 445622 194458 445706 194694
rect 445942 194458 481386 194694
rect 481622 194458 481706 194694
rect 481942 194458 517386 194694
rect 517622 194458 517706 194694
rect 517942 194458 553386 194694
rect 553622 194458 553706 194694
rect 553942 194458 588222 194694
rect 588458 194458 588542 194694
rect 588778 194458 592650 194694
rect -8726 194426 592650 194458
rect -8726 191294 592650 191326
rect -8726 191058 -3894 191294
rect -3658 191058 -3574 191294
rect -3338 191058 9666 191294
rect 9902 191058 9986 191294
rect 10222 191058 45666 191294
rect 45902 191058 45986 191294
rect 46222 191058 81666 191294
rect 81902 191058 81986 191294
rect 82222 191058 117666 191294
rect 117902 191058 117986 191294
rect 118222 191058 153666 191294
rect 153902 191058 153986 191294
rect 154222 191058 189666 191294
rect 189902 191058 189986 191294
rect 190222 191058 225666 191294
rect 225902 191058 225986 191294
rect 226222 191058 261666 191294
rect 261902 191058 261986 191294
rect 262222 191058 297666 191294
rect 297902 191058 297986 191294
rect 298222 191058 333666 191294
rect 333902 191058 333986 191294
rect 334222 191058 369666 191294
rect 369902 191058 369986 191294
rect 370222 191058 405666 191294
rect 405902 191058 405986 191294
rect 406222 191058 441666 191294
rect 441902 191058 441986 191294
rect 442222 191058 477666 191294
rect 477902 191058 477986 191294
rect 478222 191058 513666 191294
rect 513902 191058 513986 191294
rect 514222 191058 549666 191294
rect 549902 191058 549986 191294
rect 550222 191058 587262 191294
rect 587498 191058 587582 191294
rect 587818 191058 592650 191294
rect -8726 190974 592650 191058
rect -8726 190738 -3894 190974
rect -3658 190738 -3574 190974
rect -3338 190738 9666 190974
rect 9902 190738 9986 190974
rect 10222 190738 45666 190974
rect 45902 190738 45986 190974
rect 46222 190738 81666 190974
rect 81902 190738 81986 190974
rect 82222 190738 117666 190974
rect 117902 190738 117986 190974
rect 118222 190738 153666 190974
rect 153902 190738 153986 190974
rect 154222 190738 189666 190974
rect 189902 190738 189986 190974
rect 190222 190738 225666 190974
rect 225902 190738 225986 190974
rect 226222 190738 261666 190974
rect 261902 190738 261986 190974
rect 262222 190738 297666 190974
rect 297902 190738 297986 190974
rect 298222 190738 333666 190974
rect 333902 190738 333986 190974
rect 334222 190738 369666 190974
rect 369902 190738 369986 190974
rect 370222 190738 405666 190974
rect 405902 190738 405986 190974
rect 406222 190738 441666 190974
rect 441902 190738 441986 190974
rect 442222 190738 477666 190974
rect 477902 190738 477986 190974
rect 478222 190738 513666 190974
rect 513902 190738 513986 190974
rect 514222 190738 549666 190974
rect 549902 190738 549986 190974
rect 550222 190738 587262 190974
rect 587498 190738 587582 190974
rect 587818 190738 592650 190974
rect -8726 190706 592650 190738
rect -8726 187574 592650 187606
rect -8726 187338 -2934 187574
rect -2698 187338 -2614 187574
rect -2378 187338 5946 187574
rect 6182 187338 6266 187574
rect 6502 187338 41946 187574
rect 42182 187338 42266 187574
rect 42502 187338 77946 187574
rect 78182 187338 78266 187574
rect 78502 187338 99610 187574
rect 99846 187338 130330 187574
rect 130566 187338 161050 187574
rect 161286 187338 221946 187574
rect 222182 187338 222266 187574
rect 222502 187338 257946 187574
rect 258182 187338 258266 187574
rect 258502 187338 293946 187574
rect 294182 187338 294266 187574
rect 294502 187338 329946 187574
rect 330182 187338 330266 187574
rect 330502 187338 365946 187574
rect 366182 187338 366266 187574
rect 366502 187338 401946 187574
rect 402182 187338 402266 187574
rect 402502 187338 437946 187574
rect 438182 187338 438266 187574
rect 438502 187338 473946 187574
rect 474182 187338 474266 187574
rect 474502 187338 509946 187574
rect 510182 187338 510266 187574
rect 510502 187338 545946 187574
rect 546182 187338 546266 187574
rect 546502 187338 581946 187574
rect 582182 187338 582266 187574
rect 582502 187338 586302 187574
rect 586538 187338 586622 187574
rect 586858 187338 592650 187574
rect -8726 187254 592650 187338
rect -8726 187018 -2934 187254
rect -2698 187018 -2614 187254
rect -2378 187018 5946 187254
rect 6182 187018 6266 187254
rect 6502 187018 41946 187254
rect 42182 187018 42266 187254
rect 42502 187018 77946 187254
rect 78182 187018 78266 187254
rect 78502 187018 99610 187254
rect 99846 187018 130330 187254
rect 130566 187018 161050 187254
rect 161286 187018 221946 187254
rect 222182 187018 222266 187254
rect 222502 187018 257946 187254
rect 258182 187018 258266 187254
rect 258502 187018 293946 187254
rect 294182 187018 294266 187254
rect 294502 187018 329946 187254
rect 330182 187018 330266 187254
rect 330502 187018 365946 187254
rect 366182 187018 366266 187254
rect 366502 187018 401946 187254
rect 402182 187018 402266 187254
rect 402502 187018 437946 187254
rect 438182 187018 438266 187254
rect 438502 187018 473946 187254
rect 474182 187018 474266 187254
rect 474502 187018 509946 187254
rect 510182 187018 510266 187254
rect 510502 187018 545946 187254
rect 546182 187018 546266 187254
rect 546502 187018 581946 187254
rect 582182 187018 582266 187254
rect 582502 187018 586302 187254
rect 586538 187018 586622 187254
rect 586858 187018 592650 187254
rect -8726 186986 592650 187018
rect -8726 183854 592650 183886
rect -8726 183618 -1974 183854
rect -1738 183618 -1654 183854
rect -1418 183618 2226 183854
rect 2462 183618 2546 183854
rect 2782 183618 38226 183854
rect 38462 183618 38546 183854
rect 38782 183618 74226 183854
rect 74462 183618 74546 183854
rect 74782 183618 84250 183854
rect 84486 183618 114970 183854
rect 115206 183618 145690 183854
rect 145926 183618 176410 183854
rect 176646 183618 218226 183854
rect 218462 183618 218546 183854
rect 218782 183618 254226 183854
rect 254462 183618 254546 183854
rect 254782 183618 290226 183854
rect 290462 183618 290546 183854
rect 290782 183618 326226 183854
rect 326462 183618 326546 183854
rect 326782 183618 362226 183854
rect 362462 183618 362546 183854
rect 362782 183618 398226 183854
rect 398462 183618 398546 183854
rect 398782 183618 434226 183854
rect 434462 183618 434546 183854
rect 434782 183618 470226 183854
rect 470462 183618 470546 183854
rect 470782 183618 506226 183854
rect 506462 183618 506546 183854
rect 506782 183618 542226 183854
rect 542462 183618 542546 183854
rect 542782 183618 578226 183854
rect 578462 183618 578546 183854
rect 578782 183618 585342 183854
rect 585578 183618 585662 183854
rect 585898 183618 592650 183854
rect -8726 183534 592650 183618
rect -8726 183298 -1974 183534
rect -1738 183298 -1654 183534
rect -1418 183298 2226 183534
rect 2462 183298 2546 183534
rect 2782 183298 38226 183534
rect 38462 183298 38546 183534
rect 38782 183298 74226 183534
rect 74462 183298 74546 183534
rect 74782 183298 84250 183534
rect 84486 183298 114970 183534
rect 115206 183298 145690 183534
rect 145926 183298 176410 183534
rect 176646 183298 218226 183534
rect 218462 183298 218546 183534
rect 218782 183298 254226 183534
rect 254462 183298 254546 183534
rect 254782 183298 290226 183534
rect 290462 183298 290546 183534
rect 290782 183298 326226 183534
rect 326462 183298 326546 183534
rect 326782 183298 362226 183534
rect 362462 183298 362546 183534
rect 362782 183298 398226 183534
rect 398462 183298 398546 183534
rect 398782 183298 434226 183534
rect 434462 183298 434546 183534
rect 434782 183298 470226 183534
rect 470462 183298 470546 183534
rect 470782 183298 506226 183534
rect 506462 183298 506546 183534
rect 506782 183298 542226 183534
rect 542462 183298 542546 183534
rect 542782 183298 578226 183534
rect 578462 183298 578546 183534
rect 578782 183298 585342 183534
rect 585578 183298 585662 183534
rect 585898 183298 592650 183534
rect -8726 183266 592650 183298
rect -8726 173894 592650 173926
rect -8726 173658 -8694 173894
rect -8458 173658 -8374 173894
rect -8138 173658 28266 173894
rect 28502 173658 28586 173894
rect 28822 173658 64266 173894
rect 64502 173658 64586 173894
rect 64822 173658 208266 173894
rect 208502 173658 208586 173894
rect 208822 173658 244266 173894
rect 244502 173658 244586 173894
rect 244822 173658 280266 173894
rect 280502 173658 280586 173894
rect 280822 173658 316266 173894
rect 316502 173658 316586 173894
rect 316822 173658 352266 173894
rect 352502 173658 352586 173894
rect 352822 173658 388266 173894
rect 388502 173658 388586 173894
rect 388822 173658 424266 173894
rect 424502 173658 424586 173894
rect 424822 173658 460266 173894
rect 460502 173658 460586 173894
rect 460822 173658 496266 173894
rect 496502 173658 496586 173894
rect 496822 173658 532266 173894
rect 532502 173658 532586 173894
rect 532822 173658 568266 173894
rect 568502 173658 568586 173894
rect 568822 173658 592062 173894
rect 592298 173658 592382 173894
rect 592618 173658 592650 173894
rect -8726 173574 592650 173658
rect -8726 173338 -8694 173574
rect -8458 173338 -8374 173574
rect -8138 173338 28266 173574
rect 28502 173338 28586 173574
rect 28822 173338 64266 173574
rect 64502 173338 64586 173574
rect 64822 173338 208266 173574
rect 208502 173338 208586 173574
rect 208822 173338 244266 173574
rect 244502 173338 244586 173574
rect 244822 173338 280266 173574
rect 280502 173338 280586 173574
rect 280822 173338 316266 173574
rect 316502 173338 316586 173574
rect 316822 173338 352266 173574
rect 352502 173338 352586 173574
rect 352822 173338 388266 173574
rect 388502 173338 388586 173574
rect 388822 173338 424266 173574
rect 424502 173338 424586 173574
rect 424822 173338 460266 173574
rect 460502 173338 460586 173574
rect 460822 173338 496266 173574
rect 496502 173338 496586 173574
rect 496822 173338 532266 173574
rect 532502 173338 532586 173574
rect 532822 173338 568266 173574
rect 568502 173338 568586 173574
rect 568822 173338 592062 173574
rect 592298 173338 592382 173574
rect 592618 173338 592650 173574
rect -8726 173306 592650 173338
rect -8726 170174 592650 170206
rect -8726 169938 -7734 170174
rect -7498 169938 -7414 170174
rect -7178 169938 24546 170174
rect 24782 169938 24866 170174
rect 25102 169938 60546 170174
rect 60782 169938 60866 170174
rect 61102 169938 96546 170174
rect 96782 169938 96866 170174
rect 97102 169938 204546 170174
rect 204782 169938 204866 170174
rect 205102 169938 240546 170174
rect 240782 169938 240866 170174
rect 241102 169938 276546 170174
rect 276782 169938 276866 170174
rect 277102 169938 312546 170174
rect 312782 169938 312866 170174
rect 313102 169938 348546 170174
rect 348782 169938 348866 170174
rect 349102 169938 384546 170174
rect 384782 169938 384866 170174
rect 385102 169938 420546 170174
rect 420782 169938 420866 170174
rect 421102 169938 456546 170174
rect 456782 169938 456866 170174
rect 457102 169938 492546 170174
rect 492782 169938 492866 170174
rect 493102 169938 528546 170174
rect 528782 169938 528866 170174
rect 529102 169938 564546 170174
rect 564782 169938 564866 170174
rect 565102 169938 591102 170174
rect 591338 169938 591422 170174
rect 591658 169938 592650 170174
rect -8726 169854 592650 169938
rect -8726 169618 -7734 169854
rect -7498 169618 -7414 169854
rect -7178 169618 24546 169854
rect 24782 169618 24866 169854
rect 25102 169618 60546 169854
rect 60782 169618 60866 169854
rect 61102 169618 96546 169854
rect 96782 169618 96866 169854
rect 97102 169618 204546 169854
rect 204782 169618 204866 169854
rect 205102 169618 240546 169854
rect 240782 169618 240866 169854
rect 241102 169618 276546 169854
rect 276782 169618 276866 169854
rect 277102 169618 312546 169854
rect 312782 169618 312866 169854
rect 313102 169618 348546 169854
rect 348782 169618 348866 169854
rect 349102 169618 384546 169854
rect 384782 169618 384866 169854
rect 385102 169618 420546 169854
rect 420782 169618 420866 169854
rect 421102 169618 456546 169854
rect 456782 169618 456866 169854
rect 457102 169618 492546 169854
rect 492782 169618 492866 169854
rect 493102 169618 528546 169854
rect 528782 169618 528866 169854
rect 529102 169618 564546 169854
rect 564782 169618 564866 169854
rect 565102 169618 591102 169854
rect 591338 169618 591422 169854
rect 591658 169618 592650 169854
rect -8726 169586 592650 169618
rect -8726 166454 592650 166486
rect -8726 166218 -6774 166454
rect -6538 166218 -6454 166454
rect -6218 166218 20826 166454
rect 21062 166218 21146 166454
rect 21382 166218 56826 166454
rect 57062 166218 57146 166454
rect 57382 166218 92826 166454
rect 93062 166218 93146 166454
rect 93382 166218 200826 166454
rect 201062 166218 201146 166454
rect 201382 166218 236826 166454
rect 237062 166218 237146 166454
rect 237382 166218 272826 166454
rect 273062 166218 273146 166454
rect 273382 166218 308826 166454
rect 309062 166218 309146 166454
rect 309382 166218 344826 166454
rect 345062 166218 345146 166454
rect 345382 166218 380826 166454
rect 381062 166218 381146 166454
rect 381382 166218 416826 166454
rect 417062 166218 417146 166454
rect 417382 166218 452826 166454
rect 453062 166218 453146 166454
rect 453382 166218 488826 166454
rect 489062 166218 489146 166454
rect 489382 166218 524826 166454
rect 525062 166218 525146 166454
rect 525382 166218 560826 166454
rect 561062 166218 561146 166454
rect 561382 166218 590142 166454
rect 590378 166218 590462 166454
rect 590698 166218 592650 166454
rect -8726 166134 592650 166218
rect -8726 165898 -6774 166134
rect -6538 165898 -6454 166134
rect -6218 165898 20826 166134
rect 21062 165898 21146 166134
rect 21382 165898 56826 166134
rect 57062 165898 57146 166134
rect 57382 165898 92826 166134
rect 93062 165898 93146 166134
rect 93382 165898 200826 166134
rect 201062 165898 201146 166134
rect 201382 165898 236826 166134
rect 237062 165898 237146 166134
rect 237382 165898 272826 166134
rect 273062 165898 273146 166134
rect 273382 165898 308826 166134
rect 309062 165898 309146 166134
rect 309382 165898 344826 166134
rect 345062 165898 345146 166134
rect 345382 165898 380826 166134
rect 381062 165898 381146 166134
rect 381382 165898 416826 166134
rect 417062 165898 417146 166134
rect 417382 165898 452826 166134
rect 453062 165898 453146 166134
rect 453382 165898 488826 166134
rect 489062 165898 489146 166134
rect 489382 165898 524826 166134
rect 525062 165898 525146 166134
rect 525382 165898 560826 166134
rect 561062 165898 561146 166134
rect 561382 165898 590142 166134
rect 590378 165898 590462 166134
rect 590698 165898 592650 166134
rect -8726 165866 592650 165898
rect -8726 162734 592650 162766
rect -8726 162498 -5814 162734
rect -5578 162498 -5494 162734
rect -5258 162498 17106 162734
rect 17342 162498 17426 162734
rect 17662 162498 53106 162734
rect 53342 162498 53426 162734
rect 53662 162498 89106 162734
rect 89342 162498 89426 162734
rect 89662 162498 197106 162734
rect 197342 162498 197426 162734
rect 197662 162498 233106 162734
rect 233342 162498 233426 162734
rect 233662 162498 269106 162734
rect 269342 162498 269426 162734
rect 269662 162498 305106 162734
rect 305342 162498 305426 162734
rect 305662 162498 341106 162734
rect 341342 162498 341426 162734
rect 341662 162498 377106 162734
rect 377342 162498 377426 162734
rect 377662 162498 413106 162734
rect 413342 162498 413426 162734
rect 413662 162498 449106 162734
rect 449342 162498 449426 162734
rect 449662 162498 485106 162734
rect 485342 162498 485426 162734
rect 485662 162498 521106 162734
rect 521342 162498 521426 162734
rect 521662 162498 557106 162734
rect 557342 162498 557426 162734
rect 557662 162498 589182 162734
rect 589418 162498 589502 162734
rect 589738 162498 592650 162734
rect -8726 162414 592650 162498
rect -8726 162178 -5814 162414
rect -5578 162178 -5494 162414
rect -5258 162178 17106 162414
rect 17342 162178 17426 162414
rect 17662 162178 53106 162414
rect 53342 162178 53426 162414
rect 53662 162178 89106 162414
rect 89342 162178 89426 162414
rect 89662 162178 197106 162414
rect 197342 162178 197426 162414
rect 197662 162178 233106 162414
rect 233342 162178 233426 162414
rect 233662 162178 269106 162414
rect 269342 162178 269426 162414
rect 269662 162178 305106 162414
rect 305342 162178 305426 162414
rect 305662 162178 341106 162414
rect 341342 162178 341426 162414
rect 341662 162178 377106 162414
rect 377342 162178 377426 162414
rect 377662 162178 413106 162414
rect 413342 162178 413426 162414
rect 413662 162178 449106 162414
rect 449342 162178 449426 162414
rect 449662 162178 485106 162414
rect 485342 162178 485426 162414
rect 485662 162178 521106 162414
rect 521342 162178 521426 162414
rect 521662 162178 557106 162414
rect 557342 162178 557426 162414
rect 557662 162178 589182 162414
rect 589418 162178 589502 162414
rect 589738 162178 592650 162414
rect -8726 162146 592650 162178
rect -8726 159014 592650 159046
rect -8726 158778 -4854 159014
rect -4618 158778 -4534 159014
rect -4298 158778 13386 159014
rect 13622 158778 13706 159014
rect 13942 158778 49386 159014
rect 49622 158778 49706 159014
rect 49942 158778 85386 159014
rect 85622 158778 85706 159014
rect 85942 158778 193386 159014
rect 193622 158778 193706 159014
rect 193942 158778 229386 159014
rect 229622 158778 229706 159014
rect 229942 158778 265386 159014
rect 265622 158778 265706 159014
rect 265942 158778 301386 159014
rect 301622 158778 301706 159014
rect 301942 158778 337386 159014
rect 337622 158778 337706 159014
rect 337942 158778 373386 159014
rect 373622 158778 373706 159014
rect 373942 158778 409386 159014
rect 409622 158778 409706 159014
rect 409942 158778 445386 159014
rect 445622 158778 445706 159014
rect 445942 158778 481386 159014
rect 481622 158778 481706 159014
rect 481942 158778 517386 159014
rect 517622 158778 517706 159014
rect 517942 158778 553386 159014
rect 553622 158778 553706 159014
rect 553942 158778 588222 159014
rect 588458 158778 588542 159014
rect 588778 158778 592650 159014
rect -8726 158694 592650 158778
rect -8726 158458 -4854 158694
rect -4618 158458 -4534 158694
rect -4298 158458 13386 158694
rect 13622 158458 13706 158694
rect 13942 158458 49386 158694
rect 49622 158458 49706 158694
rect 49942 158458 85386 158694
rect 85622 158458 85706 158694
rect 85942 158458 193386 158694
rect 193622 158458 193706 158694
rect 193942 158458 229386 158694
rect 229622 158458 229706 158694
rect 229942 158458 265386 158694
rect 265622 158458 265706 158694
rect 265942 158458 301386 158694
rect 301622 158458 301706 158694
rect 301942 158458 337386 158694
rect 337622 158458 337706 158694
rect 337942 158458 373386 158694
rect 373622 158458 373706 158694
rect 373942 158458 409386 158694
rect 409622 158458 409706 158694
rect 409942 158458 445386 158694
rect 445622 158458 445706 158694
rect 445942 158458 481386 158694
rect 481622 158458 481706 158694
rect 481942 158458 517386 158694
rect 517622 158458 517706 158694
rect 517942 158458 553386 158694
rect 553622 158458 553706 158694
rect 553942 158458 588222 158694
rect 588458 158458 588542 158694
rect 588778 158458 592650 158694
rect -8726 158426 592650 158458
rect -8726 155294 592650 155326
rect -8726 155058 -3894 155294
rect -3658 155058 -3574 155294
rect -3338 155058 9666 155294
rect 9902 155058 9986 155294
rect 10222 155058 45666 155294
rect 45902 155058 45986 155294
rect 46222 155058 81666 155294
rect 81902 155058 81986 155294
rect 82222 155058 189666 155294
rect 189902 155058 189986 155294
rect 190222 155058 225666 155294
rect 225902 155058 225986 155294
rect 226222 155058 261666 155294
rect 261902 155058 261986 155294
rect 262222 155058 297666 155294
rect 297902 155058 297986 155294
rect 298222 155058 333666 155294
rect 333902 155058 333986 155294
rect 334222 155058 369666 155294
rect 369902 155058 369986 155294
rect 370222 155058 405666 155294
rect 405902 155058 405986 155294
rect 406222 155058 441666 155294
rect 441902 155058 441986 155294
rect 442222 155058 477666 155294
rect 477902 155058 477986 155294
rect 478222 155058 513666 155294
rect 513902 155058 513986 155294
rect 514222 155058 549666 155294
rect 549902 155058 549986 155294
rect 550222 155058 587262 155294
rect 587498 155058 587582 155294
rect 587818 155058 592650 155294
rect -8726 154974 592650 155058
rect -8726 154738 -3894 154974
rect -3658 154738 -3574 154974
rect -3338 154738 9666 154974
rect 9902 154738 9986 154974
rect 10222 154738 45666 154974
rect 45902 154738 45986 154974
rect 46222 154738 81666 154974
rect 81902 154738 81986 154974
rect 82222 154738 189666 154974
rect 189902 154738 189986 154974
rect 190222 154738 225666 154974
rect 225902 154738 225986 154974
rect 226222 154738 261666 154974
rect 261902 154738 261986 154974
rect 262222 154738 297666 154974
rect 297902 154738 297986 154974
rect 298222 154738 333666 154974
rect 333902 154738 333986 154974
rect 334222 154738 369666 154974
rect 369902 154738 369986 154974
rect 370222 154738 405666 154974
rect 405902 154738 405986 154974
rect 406222 154738 441666 154974
rect 441902 154738 441986 154974
rect 442222 154738 477666 154974
rect 477902 154738 477986 154974
rect 478222 154738 513666 154974
rect 513902 154738 513986 154974
rect 514222 154738 549666 154974
rect 549902 154738 549986 154974
rect 550222 154738 587262 154974
rect 587498 154738 587582 154974
rect 587818 154738 592650 154974
rect -8726 154706 592650 154738
rect -8726 151574 592650 151606
rect -8726 151338 -2934 151574
rect -2698 151338 -2614 151574
rect -2378 151338 5946 151574
rect 6182 151338 6266 151574
rect 6502 151338 41946 151574
rect 42182 151338 42266 151574
rect 42502 151338 77946 151574
rect 78182 151338 78266 151574
rect 78502 151338 99610 151574
rect 99846 151338 130330 151574
rect 130566 151338 161050 151574
rect 161286 151338 221946 151574
rect 222182 151338 222266 151574
rect 222502 151338 257946 151574
rect 258182 151338 258266 151574
rect 258502 151338 293946 151574
rect 294182 151338 294266 151574
rect 294502 151338 329946 151574
rect 330182 151338 330266 151574
rect 330502 151338 365946 151574
rect 366182 151338 366266 151574
rect 366502 151338 401946 151574
rect 402182 151338 402266 151574
rect 402502 151338 437946 151574
rect 438182 151338 438266 151574
rect 438502 151338 473946 151574
rect 474182 151338 474266 151574
rect 474502 151338 509946 151574
rect 510182 151338 510266 151574
rect 510502 151338 545946 151574
rect 546182 151338 546266 151574
rect 546502 151338 581946 151574
rect 582182 151338 582266 151574
rect 582502 151338 586302 151574
rect 586538 151338 586622 151574
rect 586858 151338 592650 151574
rect -8726 151254 592650 151338
rect -8726 151018 -2934 151254
rect -2698 151018 -2614 151254
rect -2378 151018 5946 151254
rect 6182 151018 6266 151254
rect 6502 151018 41946 151254
rect 42182 151018 42266 151254
rect 42502 151018 77946 151254
rect 78182 151018 78266 151254
rect 78502 151018 99610 151254
rect 99846 151018 130330 151254
rect 130566 151018 161050 151254
rect 161286 151018 221946 151254
rect 222182 151018 222266 151254
rect 222502 151018 257946 151254
rect 258182 151018 258266 151254
rect 258502 151018 293946 151254
rect 294182 151018 294266 151254
rect 294502 151018 329946 151254
rect 330182 151018 330266 151254
rect 330502 151018 365946 151254
rect 366182 151018 366266 151254
rect 366502 151018 401946 151254
rect 402182 151018 402266 151254
rect 402502 151018 437946 151254
rect 438182 151018 438266 151254
rect 438502 151018 473946 151254
rect 474182 151018 474266 151254
rect 474502 151018 509946 151254
rect 510182 151018 510266 151254
rect 510502 151018 545946 151254
rect 546182 151018 546266 151254
rect 546502 151018 581946 151254
rect 582182 151018 582266 151254
rect 582502 151018 586302 151254
rect 586538 151018 586622 151254
rect 586858 151018 592650 151254
rect -8726 150986 592650 151018
rect -8726 147854 592650 147886
rect -8726 147618 -1974 147854
rect -1738 147618 -1654 147854
rect -1418 147618 2226 147854
rect 2462 147618 2546 147854
rect 2782 147618 38226 147854
rect 38462 147618 38546 147854
rect 38782 147618 74226 147854
rect 74462 147618 74546 147854
rect 74782 147618 84250 147854
rect 84486 147618 114970 147854
rect 115206 147618 145690 147854
rect 145926 147618 176410 147854
rect 176646 147618 218226 147854
rect 218462 147618 218546 147854
rect 218782 147618 254226 147854
rect 254462 147618 254546 147854
rect 254782 147618 290226 147854
rect 290462 147618 290546 147854
rect 290782 147618 326226 147854
rect 326462 147618 326546 147854
rect 326782 147618 362226 147854
rect 362462 147618 362546 147854
rect 362782 147618 398226 147854
rect 398462 147618 398546 147854
rect 398782 147618 434226 147854
rect 434462 147618 434546 147854
rect 434782 147618 470226 147854
rect 470462 147618 470546 147854
rect 470782 147618 506226 147854
rect 506462 147618 506546 147854
rect 506782 147618 542226 147854
rect 542462 147618 542546 147854
rect 542782 147618 578226 147854
rect 578462 147618 578546 147854
rect 578782 147618 585342 147854
rect 585578 147618 585662 147854
rect 585898 147618 592650 147854
rect -8726 147534 592650 147618
rect -8726 147298 -1974 147534
rect -1738 147298 -1654 147534
rect -1418 147298 2226 147534
rect 2462 147298 2546 147534
rect 2782 147298 38226 147534
rect 38462 147298 38546 147534
rect 38782 147298 74226 147534
rect 74462 147298 74546 147534
rect 74782 147298 84250 147534
rect 84486 147298 114970 147534
rect 115206 147298 145690 147534
rect 145926 147298 176410 147534
rect 176646 147298 218226 147534
rect 218462 147298 218546 147534
rect 218782 147298 254226 147534
rect 254462 147298 254546 147534
rect 254782 147298 290226 147534
rect 290462 147298 290546 147534
rect 290782 147298 326226 147534
rect 326462 147298 326546 147534
rect 326782 147298 362226 147534
rect 362462 147298 362546 147534
rect 362782 147298 398226 147534
rect 398462 147298 398546 147534
rect 398782 147298 434226 147534
rect 434462 147298 434546 147534
rect 434782 147298 470226 147534
rect 470462 147298 470546 147534
rect 470782 147298 506226 147534
rect 506462 147298 506546 147534
rect 506782 147298 542226 147534
rect 542462 147298 542546 147534
rect 542782 147298 578226 147534
rect 578462 147298 578546 147534
rect 578782 147298 585342 147534
rect 585578 147298 585662 147534
rect 585898 147298 592650 147534
rect -8726 147266 592650 147298
rect -8726 137894 592650 137926
rect -8726 137658 -8694 137894
rect -8458 137658 -8374 137894
rect -8138 137658 28266 137894
rect 28502 137658 28586 137894
rect 28822 137658 64266 137894
rect 64502 137658 64586 137894
rect 64822 137658 208266 137894
rect 208502 137658 208586 137894
rect 208822 137658 244266 137894
rect 244502 137658 244586 137894
rect 244822 137658 280266 137894
rect 280502 137658 280586 137894
rect 280822 137658 316266 137894
rect 316502 137658 316586 137894
rect 316822 137658 352266 137894
rect 352502 137658 352586 137894
rect 352822 137658 388266 137894
rect 388502 137658 388586 137894
rect 388822 137658 424266 137894
rect 424502 137658 424586 137894
rect 424822 137658 460266 137894
rect 460502 137658 460586 137894
rect 460822 137658 496266 137894
rect 496502 137658 496586 137894
rect 496822 137658 532266 137894
rect 532502 137658 532586 137894
rect 532822 137658 568266 137894
rect 568502 137658 568586 137894
rect 568822 137658 592062 137894
rect 592298 137658 592382 137894
rect 592618 137658 592650 137894
rect -8726 137574 592650 137658
rect -8726 137338 -8694 137574
rect -8458 137338 -8374 137574
rect -8138 137338 28266 137574
rect 28502 137338 28586 137574
rect 28822 137338 64266 137574
rect 64502 137338 64586 137574
rect 64822 137338 208266 137574
rect 208502 137338 208586 137574
rect 208822 137338 244266 137574
rect 244502 137338 244586 137574
rect 244822 137338 280266 137574
rect 280502 137338 280586 137574
rect 280822 137338 316266 137574
rect 316502 137338 316586 137574
rect 316822 137338 352266 137574
rect 352502 137338 352586 137574
rect 352822 137338 388266 137574
rect 388502 137338 388586 137574
rect 388822 137338 424266 137574
rect 424502 137338 424586 137574
rect 424822 137338 460266 137574
rect 460502 137338 460586 137574
rect 460822 137338 496266 137574
rect 496502 137338 496586 137574
rect 496822 137338 532266 137574
rect 532502 137338 532586 137574
rect 532822 137338 568266 137574
rect 568502 137338 568586 137574
rect 568822 137338 592062 137574
rect 592298 137338 592382 137574
rect 592618 137338 592650 137574
rect -8726 137306 592650 137338
rect -8726 134174 592650 134206
rect -8726 133938 -7734 134174
rect -7498 133938 -7414 134174
rect -7178 133938 24546 134174
rect 24782 133938 24866 134174
rect 25102 133938 60546 134174
rect 60782 133938 60866 134174
rect 61102 133938 96546 134174
rect 96782 133938 96866 134174
rect 97102 133938 204546 134174
rect 204782 133938 204866 134174
rect 205102 133938 240546 134174
rect 240782 133938 240866 134174
rect 241102 133938 276546 134174
rect 276782 133938 276866 134174
rect 277102 133938 312546 134174
rect 312782 133938 312866 134174
rect 313102 133938 348546 134174
rect 348782 133938 348866 134174
rect 349102 133938 384546 134174
rect 384782 133938 384866 134174
rect 385102 133938 420546 134174
rect 420782 133938 420866 134174
rect 421102 133938 456546 134174
rect 456782 133938 456866 134174
rect 457102 133938 492546 134174
rect 492782 133938 492866 134174
rect 493102 133938 528546 134174
rect 528782 133938 528866 134174
rect 529102 133938 564546 134174
rect 564782 133938 564866 134174
rect 565102 133938 591102 134174
rect 591338 133938 591422 134174
rect 591658 133938 592650 134174
rect -8726 133854 592650 133938
rect -8726 133618 -7734 133854
rect -7498 133618 -7414 133854
rect -7178 133618 24546 133854
rect 24782 133618 24866 133854
rect 25102 133618 60546 133854
rect 60782 133618 60866 133854
rect 61102 133618 96546 133854
rect 96782 133618 96866 133854
rect 97102 133618 204546 133854
rect 204782 133618 204866 133854
rect 205102 133618 240546 133854
rect 240782 133618 240866 133854
rect 241102 133618 276546 133854
rect 276782 133618 276866 133854
rect 277102 133618 312546 133854
rect 312782 133618 312866 133854
rect 313102 133618 348546 133854
rect 348782 133618 348866 133854
rect 349102 133618 384546 133854
rect 384782 133618 384866 133854
rect 385102 133618 420546 133854
rect 420782 133618 420866 133854
rect 421102 133618 456546 133854
rect 456782 133618 456866 133854
rect 457102 133618 492546 133854
rect 492782 133618 492866 133854
rect 493102 133618 528546 133854
rect 528782 133618 528866 133854
rect 529102 133618 564546 133854
rect 564782 133618 564866 133854
rect 565102 133618 591102 133854
rect 591338 133618 591422 133854
rect 591658 133618 592650 133854
rect -8726 133586 592650 133618
rect -8726 130454 592650 130486
rect -8726 130218 -6774 130454
rect -6538 130218 -6454 130454
rect -6218 130218 20826 130454
rect 21062 130218 21146 130454
rect 21382 130218 56826 130454
rect 57062 130218 57146 130454
rect 57382 130218 92826 130454
rect 93062 130218 93146 130454
rect 93382 130218 200826 130454
rect 201062 130218 201146 130454
rect 201382 130218 236826 130454
rect 237062 130218 237146 130454
rect 237382 130218 272826 130454
rect 273062 130218 273146 130454
rect 273382 130218 308826 130454
rect 309062 130218 309146 130454
rect 309382 130218 344826 130454
rect 345062 130218 345146 130454
rect 345382 130218 380826 130454
rect 381062 130218 381146 130454
rect 381382 130218 452826 130454
rect 453062 130218 453146 130454
rect 453382 130218 488826 130454
rect 489062 130218 489146 130454
rect 489382 130218 524826 130454
rect 525062 130218 525146 130454
rect 525382 130218 560826 130454
rect 561062 130218 561146 130454
rect 561382 130218 590142 130454
rect 590378 130218 590462 130454
rect 590698 130218 592650 130454
rect -8726 130134 592650 130218
rect -8726 129898 -6774 130134
rect -6538 129898 -6454 130134
rect -6218 129898 20826 130134
rect 21062 129898 21146 130134
rect 21382 129898 56826 130134
rect 57062 129898 57146 130134
rect 57382 129898 92826 130134
rect 93062 129898 93146 130134
rect 93382 129898 200826 130134
rect 201062 129898 201146 130134
rect 201382 129898 236826 130134
rect 237062 129898 237146 130134
rect 237382 129898 272826 130134
rect 273062 129898 273146 130134
rect 273382 129898 308826 130134
rect 309062 129898 309146 130134
rect 309382 129898 344826 130134
rect 345062 129898 345146 130134
rect 345382 129898 380826 130134
rect 381062 129898 381146 130134
rect 381382 129898 452826 130134
rect 453062 129898 453146 130134
rect 453382 129898 488826 130134
rect 489062 129898 489146 130134
rect 489382 129898 524826 130134
rect 525062 129898 525146 130134
rect 525382 129898 560826 130134
rect 561062 129898 561146 130134
rect 561382 129898 590142 130134
rect 590378 129898 590462 130134
rect 590698 129898 592650 130134
rect -8726 129866 592650 129898
rect -8726 126734 592650 126766
rect -8726 126498 -5814 126734
rect -5578 126498 -5494 126734
rect -5258 126498 17106 126734
rect 17342 126498 17426 126734
rect 17662 126498 53106 126734
rect 53342 126498 53426 126734
rect 53662 126498 89106 126734
rect 89342 126498 89426 126734
rect 89662 126498 197106 126734
rect 197342 126498 197426 126734
rect 197662 126498 233106 126734
rect 233342 126498 233426 126734
rect 233662 126498 269106 126734
rect 269342 126498 269426 126734
rect 269662 126498 305106 126734
rect 305342 126498 305426 126734
rect 305662 126498 341106 126734
rect 341342 126498 341426 126734
rect 341662 126498 377106 126734
rect 377342 126498 377426 126734
rect 377662 126498 485106 126734
rect 485342 126498 485426 126734
rect 485662 126498 521106 126734
rect 521342 126498 521426 126734
rect 521662 126498 557106 126734
rect 557342 126498 557426 126734
rect 557662 126498 589182 126734
rect 589418 126498 589502 126734
rect 589738 126498 592650 126734
rect -8726 126414 592650 126498
rect -8726 126178 -5814 126414
rect -5578 126178 -5494 126414
rect -5258 126178 17106 126414
rect 17342 126178 17426 126414
rect 17662 126178 53106 126414
rect 53342 126178 53426 126414
rect 53662 126178 89106 126414
rect 89342 126178 89426 126414
rect 89662 126178 197106 126414
rect 197342 126178 197426 126414
rect 197662 126178 233106 126414
rect 233342 126178 233426 126414
rect 233662 126178 269106 126414
rect 269342 126178 269426 126414
rect 269662 126178 305106 126414
rect 305342 126178 305426 126414
rect 305662 126178 341106 126414
rect 341342 126178 341426 126414
rect 341662 126178 377106 126414
rect 377342 126178 377426 126414
rect 377662 126178 485106 126414
rect 485342 126178 485426 126414
rect 485662 126178 521106 126414
rect 521342 126178 521426 126414
rect 521662 126178 557106 126414
rect 557342 126178 557426 126414
rect 557662 126178 589182 126414
rect 589418 126178 589502 126414
rect 589738 126178 592650 126414
rect -8726 126146 592650 126178
rect -8726 123014 592650 123046
rect -8726 122778 -4854 123014
rect -4618 122778 -4534 123014
rect -4298 122778 13386 123014
rect 13622 122778 13706 123014
rect 13942 122778 49386 123014
rect 49622 122778 49706 123014
rect 49942 122778 85386 123014
rect 85622 122778 85706 123014
rect 85942 122778 193386 123014
rect 193622 122778 193706 123014
rect 193942 122778 229386 123014
rect 229622 122778 229706 123014
rect 229942 122778 265386 123014
rect 265622 122778 265706 123014
rect 265942 122778 301386 123014
rect 301622 122778 301706 123014
rect 301942 122778 337386 123014
rect 337622 122778 337706 123014
rect 337942 122778 373386 123014
rect 373622 122778 373706 123014
rect 373942 122778 409386 123014
rect 409622 122778 409706 123014
rect 409942 122778 481386 123014
rect 481622 122778 481706 123014
rect 481942 122778 517386 123014
rect 517622 122778 517706 123014
rect 517942 122778 553386 123014
rect 553622 122778 553706 123014
rect 553942 122778 588222 123014
rect 588458 122778 588542 123014
rect 588778 122778 592650 123014
rect -8726 122694 592650 122778
rect -8726 122458 -4854 122694
rect -4618 122458 -4534 122694
rect -4298 122458 13386 122694
rect 13622 122458 13706 122694
rect 13942 122458 49386 122694
rect 49622 122458 49706 122694
rect 49942 122458 85386 122694
rect 85622 122458 85706 122694
rect 85942 122458 193386 122694
rect 193622 122458 193706 122694
rect 193942 122458 229386 122694
rect 229622 122458 229706 122694
rect 229942 122458 265386 122694
rect 265622 122458 265706 122694
rect 265942 122458 301386 122694
rect 301622 122458 301706 122694
rect 301942 122458 337386 122694
rect 337622 122458 337706 122694
rect 337942 122458 373386 122694
rect 373622 122458 373706 122694
rect 373942 122458 409386 122694
rect 409622 122458 409706 122694
rect 409942 122458 481386 122694
rect 481622 122458 481706 122694
rect 481942 122458 517386 122694
rect 517622 122458 517706 122694
rect 517942 122458 553386 122694
rect 553622 122458 553706 122694
rect 553942 122458 588222 122694
rect 588458 122458 588542 122694
rect 588778 122458 592650 122694
rect -8726 122426 592650 122458
rect -8726 119294 592650 119326
rect -8726 119058 -3894 119294
rect -3658 119058 -3574 119294
rect -3338 119058 9666 119294
rect 9902 119058 9986 119294
rect 10222 119058 45666 119294
rect 45902 119058 45986 119294
rect 46222 119058 81666 119294
rect 81902 119058 81986 119294
rect 82222 119058 189666 119294
rect 189902 119058 189986 119294
rect 190222 119058 225666 119294
rect 225902 119058 225986 119294
rect 226222 119058 261666 119294
rect 261902 119058 261986 119294
rect 262222 119058 297666 119294
rect 297902 119058 297986 119294
rect 298222 119058 333666 119294
rect 333902 119058 333986 119294
rect 334222 119058 369666 119294
rect 369902 119058 369986 119294
rect 370222 119058 405666 119294
rect 405902 119058 405986 119294
rect 406222 119058 477666 119294
rect 477902 119058 477986 119294
rect 478222 119058 513666 119294
rect 513902 119058 513986 119294
rect 514222 119058 549666 119294
rect 549902 119058 549986 119294
rect 550222 119058 587262 119294
rect 587498 119058 587582 119294
rect 587818 119058 592650 119294
rect -8726 118974 592650 119058
rect -8726 118738 -3894 118974
rect -3658 118738 -3574 118974
rect -3338 118738 9666 118974
rect 9902 118738 9986 118974
rect 10222 118738 45666 118974
rect 45902 118738 45986 118974
rect 46222 118738 81666 118974
rect 81902 118738 81986 118974
rect 82222 118738 189666 118974
rect 189902 118738 189986 118974
rect 190222 118738 225666 118974
rect 225902 118738 225986 118974
rect 226222 118738 261666 118974
rect 261902 118738 261986 118974
rect 262222 118738 297666 118974
rect 297902 118738 297986 118974
rect 298222 118738 333666 118974
rect 333902 118738 333986 118974
rect 334222 118738 369666 118974
rect 369902 118738 369986 118974
rect 370222 118738 405666 118974
rect 405902 118738 405986 118974
rect 406222 118738 477666 118974
rect 477902 118738 477986 118974
rect 478222 118738 513666 118974
rect 513902 118738 513986 118974
rect 514222 118738 549666 118974
rect 549902 118738 549986 118974
rect 550222 118738 587262 118974
rect 587498 118738 587582 118974
rect 587818 118738 592650 118974
rect -8726 118706 592650 118738
rect -8726 115574 592650 115606
rect -8726 115338 -2934 115574
rect -2698 115338 -2614 115574
rect -2378 115338 5946 115574
rect 6182 115338 6266 115574
rect 6502 115338 41946 115574
rect 42182 115338 42266 115574
rect 42502 115338 77946 115574
rect 78182 115338 78266 115574
rect 78502 115338 99610 115574
rect 99846 115338 130330 115574
rect 130566 115338 161050 115574
rect 161286 115338 221946 115574
rect 222182 115338 222266 115574
rect 222502 115338 257946 115574
rect 258182 115338 258266 115574
rect 258502 115338 293946 115574
rect 294182 115338 294266 115574
rect 294502 115338 319610 115574
rect 319846 115338 329946 115574
rect 330182 115338 330266 115574
rect 330502 115338 365946 115574
rect 366182 115338 366266 115574
rect 366502 115338 401946 115574
rect 402182 115338 402266 115574
rect 402502 115338 419610 115574
rect 419846 115338 450330 115574
rect 450566 115338 473946 115574
rect 474182 115338 474266 115574
rect 474502 115338 509946 115574
rect 510182 115338 510266 115574
rect 510502 115338 545946 115574
rect 546182 115338 546266 115574
rect 546502 115338 581946 115574
rect 582182 115338 582266 115574
rect 582502 115338 586302 115574
rect 586538 115338 586622 115574
rect 586858 115338 592650 115574
rect -8726 115254 592650 115338
rect -8726 115018 -2934 115254
rect -2698 115018 -2614 115254
rect -2378 115018 5946 115254
rect 6182 115018 6266 115254
rect 6502 115018 41946 115254
rect 42182 115018 42266 115254
rect 42502 115018 77946 115254
rect 78182 115018 78266 115254
rect 78502 115018 99610 115254
rect 99846 115018 130330 115254
rect 130566 115018 161050 115254
rect 161286 115018 221946 115254
rect 222182 115018 222266 115254
rect 222502 115018 257946 115254
rect 258182 115018 258266 115254
rect 258502 115018 293946 115254
rect 294182 115018 294266 115254
rect 294502 115018 319610 115254
rect 319846 115018 329946 115254
rect 330182 115018 330266 115254
rect 330502 115018 365946 115254
rect 366182 115018 366266 115254
rect 366502 115018 401946 115254
rect 402182 115018 402266 115254
rect 402502 115018 419610 115254
rect 419846 115018 450330 115254
rect 450566 115018 473946 115254
rect 474182 115018 474266 115254
rect 474502 115018 509946 115254
rect 510182 115018 510266 115254
rect 510502 115018 545946 115254
rect 546182 115018 546266 115254
rect 546502 115018 581946 115254
rect 582182 115018 582266 115254
rect 582502 115018 586302 115254
rect 586538 115018 586622 115254
rect 586858 115018 592650 115254
rect -8726 114986 592650 115018
rect -8726 111854 592650 111886
rect -8726 111618 -1974 111854
rect -1738 111618 -1654 111854
rect -1418 111618 2226 111854
rect 2462 111618 2546 111854
rect 2782 111618 38226 111854
rect 38462 111618 38546 111854
rect 38782 111618 74226 111854
rect 74462 111618 74546 111854
rect 74782 111618 84250 111854
rect 84486 111618 114970 111854
rect 115206 111618 145690 111854
rect 145926 111618 176410 111854
rect 176646 111618 218226 111854
rect 218462 111618 218546 111854
rect 218782 111618 254226 111854
rect 254462 111618 254546 111854
rect 254782 111618 290226 111854
rect 290462 111618 290546 111854
rect 290782 111618 304250 111854
rect 304486 111618 326226 111854
rect 326462 111618 326546 111854
rect 326782 111618 334970 111854
rect 335206 111618 362226 111854
rect 362462 111618 362546 111854
rect 362782 111618 398226 111854
rect 398462 111618 398546 111854
rect 398782 111618 404250 111854
rect 404486 111618 434970 111854
rect 435206 111618 470226 111854
rect 470462 111618 470546 111854
rect 470782 111618 506226 111854
rect 506462 111618 506546 111854
rect 506782 111618 542226 111854
rect 542462 111618 542546 111854
rect 542782 111618 578226 111854
rect 578462 111618 578546 111854
rect 578782 111618 585342 111854
rect 585578 111618 585662 111854
rect 585898 111618 592650 111854
rect -8726 111534 592650 111618
rect -8726 111298 -1974 111534
rect -1738 111298 -1654 111534
rect -1418 111298 2226 111534
rect 2462 111298 2546 111534
rect 2782 111298 38226 111534
rect 38462 111298 38546 111534
rect 38782 111298 74226 111534
rect 74462 111298 74546 111534
rect 74782 111298 84250 111534
rect 84486 111298 114970 111534
rect 115206 111298 145690 111534
rect 145926 111298 176410 111534
rect 176646 111298 218226 111534
rect 218462 111298 218546 111534
rect 218782 111298 254226 111534
rect 254462 111298 254546 111534
rect 254782 111298 290226 111534
rect 290462 111298 290546 111534
rect 290782 111298 304250 111534
rect 304486 111298 326226 111534
rect 326462 111298 326546 111534
rect 326782 111298 334970 111534
rect 335206 111298 362226 111534
rect 362462 111298 362546 111534
rect 362782 111298 398226 111534
rect 398462 111298 398546 111534
rect 398782 111298 404250 111534
rect 404486 111298 434970 111534
rect 435206 111298 470226 111534
rect 470462 111298 470546 111534
rect 470782 111298 506226 111534
rect 506462 111298 506546 111534
rect 506782 111298 542226 111534
rect 542462 111298 542546 111534
rect 542782 111298 578226 111534
rect 578462 111298 578546 111534
rect 578782 111298 585342 111534
rect 585578 111298 585662 111534
rect 585898 111298 592650 111534
rect -8726 111266 592650 111298
rect -8726 101894 592650 101926
rect -8726 101658 -8694 101894
rect -8458 101658 -8374 101894
rect -8138 101658 28266 101894
rect 28502 101658 28586 101894
rect 28822 101658 64266 101894
rect 64502 101658 64586 101894
rect 64822 101658 208266 101894
rect 208502 101658 208586 101894
rect 208822 101658 244266 101894
rect 244502 101658 244586 101894
rect 244822 101658 280266 101894
rect 280502 101658 280586 101894
rect 280822 101658 316266 101894
rect 316502 101658 316586 101894
rect 316822 101658 352266 101894
rect 352502 101658 352586 101894
rect 352822 101658 388266 101894
rect 388502 101658 388586 101894
rect 388822 101658 460266 101894
rect 460502 101658 460586 101894
rect 460822 101658 496266 101894
rect 496502 101658 496586 101894
rect 496822 101658 532266 101894
rect 532502 101658 532586 101894
rect 532822 101658 568266 101894
rect 568502 101658 568586 101894
rect 568822 101658 592062 101894
rect 592298 101658 592382 101894
rect 592618 101658 592650 101894
rect -8726 101574 592650 101658
rect -8726 101338 -8694 101574
rect -8458 101338 -8374 101574
rect -8138 101338 28266 101574
rect 28502 101338 28586 101574
rect 28822 101338 64266 101574
rect 64502 101338 64586 101574
rect 64822 101338 208266 101574
rect 208502 101338 208586 101574
rect 208822 101338 244266 101574
rect 244502 101338 244586 101574
rect 244822 101338 280266 101574
rect 280502 101338 280586 101574
rect 280822 101338 316266 101574
rect 316502 101338 316586 101574
rect 316822 101338 352266 101574
rect 352502 101338 352586 101574
rect 352822 101338 388266 101574
rect 388502 101338 388586 101574
rect 388822 101338 460266 101574
rect 460502 101338 460586 101574
rect 460822 101338 496266 101574
rect 496502 101338 496586 101574
rect 496822 101338 532266 101574
rect 532502 101338 532586 101574
rect 532822 101338 568266 101574
rect 568502 101338 568586 101574
rect 568822 101338 592062 101574
rect 592298 101338 592382 101574
rect 592618 101338 592650 101574
rect -8726 101306 592650 101338
rect -8726 98174 592650 98206
rect -8726 97938 -7734 98174
rect -7498 97938 -7414 98174
rect -7178 97938 24546 98174
rect 24782 97938 24866 98174
rect 25102 97938 60546 98174
rect 60782 97938 60866 98174
rect 61102 97938 96546 98174
rect 96782 97938 96866 98174
rect 97102 97938 204546 98174
rect 204782 97938 204866 98174
rect 205102 97938 240546 98174
rect 240782 97938 240866 98174
rect 241102 97938 276546 98174
rect 276782 97938 276866 98174
rect 277102 97938 312546 98174
rect 312782 97938 312866 98174
rect 313102 97938 348546 98174
rect 348782 97938 348866 98174
rect 349102 97938 384546 98174
rect 384782 97938 384866 98174
rect 385102 97938 456546 98174
rect 456782 97938 456866 98174
rect 457102 97938 492546 98174
rect 492782 97938 492866 98174
rect 493102 97938 528546 98174
rect 528782 97938 528866 98174
rect 529102 97938 564546 98174
rect 564782 97938 564866 98174
rect 565102 97938 591102 98174
rect 591338 97938 591422 98174
rect 591658 97938 592650 98174
rect -8726 97854 592650 97938
rect -8726 97618 -7734 97854
rect -7498 97618 -7414 97854
rect -7178 97618 24546 97854
rect 24782 97618 24866 97854
rect 25102 97618 60546 97854
rect 60782 97618 60866 97854
rect 61102 97618 96546 97854
rect 96782 97618 96866 97854
rect 97102 97618 204546 97854
rect 204782 97618 204866 97854
rect 205102 97618 240546 97854
rect 240782 97618 240866 97854
rect 241102 97618 276546 97854
rect 276782 97618 276866 97854
rect 277102 97618 312546 97854
rect 312782 97618 312866 97854
rect 313102 97618 348546 97854
rect 348782 97618 348866 97854
rect 349102 97618 384546 97854
rect 384782 97618 384866 97854
rect 385102 97618 456546 97854
rect 456782 97618 456866 97854
rect 457102 97618 492546 97854
rect 492782 97618 492866 97854
rect 493102 97618 528546 97854
rect 528782 97618 528866 97854
rect 529102 97618 564546 97854
rect 564782 97618 564866 97854
rect 565102 97618 591102 97854
rect 591338 97618 591422 97854
rect 591658 97618 592650 97854
rect -8726 97586 592650 97618
rect -8726 94454 592650 94486
rect -8726 94218 -6774 94454
rect -6538 94218 -6454 94454
rect -6218 94218 20826 94454
rect 21062 94218 21146 94454
rect 21382 94218 56826 94454
rect 57062 94218 57146 94454
rect 57382 94218 92826 94454
rect 93062 94218 93146 94454
rect 93382 94218 200826 94454
rect 201062 94218 201146 94454
rect 201382 94218 236826 94454
rect 237062 94218 237146 94454
rect 237382 94218 272826 94454
rect 273062 94218 273146 94454
rect 273382 94218 308826 94454
rect 309062 94218 309146 94454
rect 309382 94218 344826 94454
rect 345062 94218 345146 94454
rect 345382 94218 380826 94454
rect 381062 94218 381146 94454
rect 381382 94218 452826 94454
rect 453062 94218 453146 94454
rect 453382 94218 488826 94454
rect 489062 94218 489146 94454
rect 489382 94218 524826 94454
rect 525062 94218 525146 94454
rect 525382 94218 560826 94454
rect 561062 94218 561146 94454
rect 561382 94218 590142 94454
rect 590378 94218 590462 94454
rect 590698 94218 592650 94454
rect -8726 94134 592650 94218
rect -8726 93898 -6774 94134
rect -6538 93898 -6454 94134
rect -6218 93898 20826 94134
rect 21062 93898 21146 94134
rect 21382 93898 56826 94134
rect 57062 93898 57146 94134
rect 57382 93898 92826 94134
rect 93062 93898 93146 94134
rect 93382 93898 200826 94134
rect 201062 93898 201146 94134
rect 201382 93898 236826 94134
rect 237062 93898 237146 94134
rect 237382 93898 272826 94134
rect 273062 93898 273146 94134
rect 273382 93898 308826 94134
rect 309062 93898 309146 94134
rect 309382 93898 344826 94134
rect 345062 93898 345146 94134
rect 345382 93898 380826 94134
rect 381062 93898 381146 94134
rect 381382 93898 452826 94134
rect 453062 93898 453146 94134
rect 453382 93898 488826 94134
rect 489062 93898 489146 94134
rect 489382 93898 524826 94134
rect 525062 93898 525146 94134
rect 525382 93898 560826 94134
rect 561062 93898 561146 94134
rect 561382 93898 590142 94134
rect 590378 93898 590462 94134
rect 590698 93898 592650 94134
rect -8726 93866 592650 93898
rect -8726 90734 592650 90766
rect -8726 90498 -5814 90734
rect -5578 90498 -5494 90734
rect -5258 90498 17106 90734
rect 17342 90498 17426 90734
rect 17662 90498 53106 90734
rect 53342 90498 53426 90734
rect 53662 90498 89106 90734
rect 89342 90498 89426 90734
rect 89662 90498 197106 90734
rect 197342 90498 197426 90734
rect 197662 90498 233106 90734
rect 233342 90498 233426 90734
rect 233662 90498 269106 90734
rect 269342 90498 269426 90734
rect 269662 90498 305106 90734
rect 305342 90498 305426 90734
rect 305662 90498 341106 90734
rect 341342 90498 341426 90734
rect 341662 90498 377106 90734
rect 377342 90498 377426 90734
rect 377662 90498 485106 90734
rect 485342 90498 485426 90734
rect 485662 90498 521106 90734
rect 521342 90498 521426 90734
rect 521662 90498 557106 90734
rect 557342 90498 557426 90734
rect 557662 90498 589182 90734
rect 589418 90498 589502 90734
rect 589738 90498 592650 90734
rect -8726 90414 592650 90498
rect -8726 90178 -5814 90414
rect -5578 90178 -5494 90414
rect -5258 90178 17106 90414
rect 17342 90178 17426 90414
rect 17662 90178 53106 90414
rect 53342 90178 53426 90414
rect 53662 90178 89106 90414
rect 89342 90178 89426 90414
rect 89662 90178 197106 90414
rect 197342 90178 197426 90414
rect 197662 90178 233106 90414
rect 233342 90178 233426 90414
rect 233662 90178 269106 90414
rect 269342 90178 269426 90414
rect 269662 90178 305106 90414
rect 305342 90178 305426 90414
rect 305662 90178 341106 90414
rect 341342 90178 341426 90414
rect 341662 90178 377106 90414
rect 377342 90178 377426 90414
rect 377662 90178 485106 90414
rect 485342 90178 485426 90414
rect 485662 90178 521106 90414
rect 521342 90178 521426 90414
rect 521662 90178 557106 90414
rect 557342 90178 557426 90414
rect 557662 90178 589182 90414
rect 589418 90178 589502 90414
rect 589738 90178 592650 90414
rect -8726 90146 592650 90178
rect -8726 87014 592650 87046
rect -8726 86778 -4854 87014
rect -4618 86778 -4534 87014
rect -4298 86778 13386 87014
rect 13622 86778 13706 87014
rect 13942 86778 49386 87014
rect 49622 86778 49706 87014
rect 49942 86778 85386 87014
rect 85622 86778 85706 87014
rect 85942 86778 193386 87014
rect 193622 86778 193706 87014
rect 193942 86778 229386 87014
rect 229622 86778 229706 87014
rect 229942 86778 265386 87014
rect 265622 86778 265706 87014
rect 265942 86778 301386 87014
rect 301622 86778 301706 87014
rect 301942 86778 337386 87014
rect 337622 86778 337706 87014
rect 337942 86778 373386 87014
rect 373622 86778 373706 87014
rect 373942 86778 409386 87014
rect 409622 86778 409706 87014
rect 409942 86778 481386 87014
rect 481622 86778 481706 87014
rect 481942 86778 517386 87014
rect 517622 86778 517706 87014
rect 517942 86778 553386 87014
rect 553622 86778 553706 87014
rect 553942 86778 588222 87014
rect 588458 86778 588542 87014
rect 588778 86778 592650 87014
rect -8726 86694 592650 86778
rect -8726 86458 -4854 86694
rect -4618 86458 -4534 86694
rect -4298 86458 13386 86694
rect 13622 86458 13706 86694
rect 13942 86458 49386 86694
rect 49622 86458 49706 86694
rect 49942 86458 85386 86694
rect 85622 86458 85706 86694
rect 85942 86458 193386 86694
rect 193622 86458 193706 86694
rect 193942 86458 229386 86694
rect 229622 86458 229706 86694
rect 229942 86458 265386 86694
rect 265622 86458 265706 86694
rect 265942 86458 301386 86694
rect 301622 86458 301706 86694
rect 301942 86458 337386 86694
rect 337622 86458 337706 86694
rect 337942 86458 373386 86694
rect 373622 86458 373706 86694
rect 373942 86458 409386 86694
rect 409622 86458 409706 86694
rect 409942 86458 481386 86694
rect 481622 86458 481706 86694
rect 481942 86458 517386 86694
rect 517622 86458 517706 86694
rect 517942 86458 553386 86694
rect 553622 86458 553706 86694
rect 553942 86458 588222 86694
rect 588458 86458 588542 86694
rect 588778 86458 592650 86694
rect -8726 86426 592650 86458
rect -8726 83294 592650 83326
rect -8726 83058 -3894 83294
rect -3658 83058 -3574 83294
rect -3338 83058 9666 83294
rect 9902 83058 9986 83294
rect 10222 83058 45666 83294
rect 45902 83058 45986 83294
rect 46222 83058 81666 83294
rect 81902 83058 81986 83294
rect 82222 83058 189666 83294
rect 189902 83058 189986 83294
rect 190222 83058 225666 83294
rect 225902 83058 225986 83294
rect 226222 83058 261666 83294
rect 261902 83058 261986 83294
rect 262222 83058 297666 83294
rect 297902 83058 297986 83294
rect 298222 83058 333666 83294
rect 333902 83058 333986 83294
rect 334222 83058 369666 83294
rect 369902 83058 369986 83294
rect 370222 83058 405666 83294
rect 405902 83058 405986 83294
rect 406222 83058 477666 83294
rect 477902 83058 477986 83294
rect 478222 83058 513666 83294
rect 513902 83058 513986 83294
rect 514222 83058 549666 83294
rect 549902 83058 549986 83294
rect 550222 83058 587262 83294
rect 587498 83058 587582 83294
rect 587818 83058 592650 83294
rect -8726 82974 592650 83058
rect -8726 82738 -3894 82974
rect -3658 82738 -3574 82974
rect -3338 82738 9666 82974
rect 9902 82738 9986 82974
rect 10222 82738 45666 82974
rect 45902 82738 45986 82974
rect 46222 82738 81666 82974
rect 81902 82738 81986 82974
rect 82222 82738 189666 82974
rect 189902 82738 189986 82974
rect 190222 82738 225666 82974
rect 225902 82738 225986 82974
rect 226222 82738 261666 82974
rect 261902 82738 261986 82974
rect 262222 82738 297666 82974
rect 297902 82738 297986 82974
rect 298222 82738 333666 82974
rect 333902 82738 333986 82974
rect 334222 82738 369666 82974
rect 369902 82738 369986 82974
rect 370222 82738 405666 82974
rect 405902 82738 405986 82974
rect 406222 82738 477666 82974
rect 477902 82738 477986 82974
rect 478222 82738 513666 82974
rect 513902 82738 513986 82974
rect 514222 82738 549666 82974
rect 549902 82738 549986 82974
rect 550222 82738 587262 82974
rect 587498 82738 587582 82974
rect 587818 82738 592650 82974
rect -8726 82706 592650 82738
rect -8726 79574 592650 79606
rect -8726 79338 -2934 79574
rect -2698 79338 -2614 79574
rect -2378 79338 5946 79574
rect 6182 79338 6266 79574
rect 6502 79338 41946 79574
rect 42182 79338 42266 79574
rect 42502 79338 77946 79574
rect 78182 79338 78266 79574
rect 78502 79338 113946 79574
rect 114182 79338 114266 79574
rect 114502 79338 149946 79574
rect 150182 79338 150266 79574
rect 150502 79338 185946 79574
rect 186182 79338 186266 79574
rect 186502 79338 221946 79574
rect 222182 79338 222266 79574
rect 222502 79338 257946 79574
rect 258182 79338 258266 79574
rect 258502 79338 293946 79574
rect 294182 79338 294266 79574
rect 294502 79338 329946 79574
rect 330182 79338 330266 79574
rect 330502 79338 365946 79574
rect 366182 79338 366266 79574
rect 366502 79338 401946 79574
rect 402182 79338 402266 79574
rect 402502 79338 437946 79574
rect 438182 79338 438266 79574
rect 438502 79338 473946 79574
rect 474182 79338 474266 79574
rect 474502 79338 509946 79574
rect 510182 79338 510266 79574
rect 510502 79338 545946 79574
rect 546182 79338 546266 79574
rect 546502 79338 581946 79574
rect 582182 79338 582266 79574
rect 582502 79338 586302 79574
rect 586538 79338 586622 79574
rect 586858 79338 592650 79574
rect -8726 79254 592650 79338
rect -8726 79018 -2934 79254
rect -2698 79018 -2614 79254
rect -2378 79018 5946 79254
rect 6182 79018 6266 79254
rect 6502 79018 41946 79254
rect 42182 79018 42266 79254
rect 42502 79018 77946 79254
rect 78182 79018 78266 79254
rect 78502 79018 113946 79254
rect 114182 79018 114266 79254
rect 114502 79018 149946 79254
rect 150182 79018 150266 79254
rect 150502 79018 185946 79254
rect 186182 79018 186266 79254
rect 186502 79018 221946 79254
rect 222182 79018 222266 79254
rect 222502 79018 257946 79254
rect 258182 79018 258266 79254
rect 258502 79018 293946 79254
rect 294182 79018 294266 79254
rect 294502 79018 329946 79254
rect 330182 79018 330266 79254
rect 330502 79018 365946 79254
rect 366182 79018 366266 79254
rect 366502 79018 401946 79254
rect 402182 79018 402266 79254
rect 402502 79018 437946 79254
rect 438182 79018 438266 79254
rect 438502 79018 473946 79254
rect 474182 79018 474266 79254
rect 474502 79018 509946 79254
rect 510182 79018 510266 79254
rect 510502 79018 545946 79254
rect 546182 79018 546266 79254
rect 546502 79018 581946 79254
rect 582182 79018 582266 79254
rect 582502 79018 586302 79254
rect 586538 79018 586622 79254
rect 586858 79018 592650 79254
rect -8726 78986 592650 79018
rect 94876 77978 175420 78020
rect 94876 77742 94918 77978
rect 95154 77742 175142 77978
rect 175378 77742 175420 77978
rect 94876 77700 175420 77742
rect 177124 77978 324460 78020
rect 177124 77742 177166 77978
rect 177402 77742 324182 77978
rect 324418 77742 324460 77978
rect 177124 77700 324460 77742
rect -8726 75854 592650 75886
rect -8726 75618 -1974 75854
rect -1738 75618 -1654 75854
rect -1418 75618 2226 75854
rect 2462 75618 2546 75854
rect 2782 75618 38226 75854
rect 38462 75618 38546 75854
rect 38782 75618 74226 75854
rect 74462 75618 74546 75854
rect 74782 75618 110226 75854
rect 110462 75618 110546 75854
rect 110782 75618 146226 75854
rect 146462 75618 146546 75854
rect 146782 75618 182226 75854
rect 182462 75618 182546 75854
rect 182782 75618 218226 75854
rect 218462 75618 218546 75854
rect 218782 75618 254226 75854
rect 254462 75618 254546 75854
rect 254782 75618 290226 75854
rect 290462 75618 290546 75854
rect 290782 75618 326226 75854
rect 326462 75618 326546 75854
rect 326782 75618 362226 75854
rect 362462 75618 362546 75854
rect 362782 75618 398226 75854
rect 398462 75618 398546 75854
rect 398782 75618 434226 75854
rect 434462 75618 434546 75854
rect 434782 75618 470226 75854
rect 470462 75618 470546 75854
rect 470782 75618 506226 75854
rect 506462 75618 506546 75854
rect 506782 75618 542226 75854
rect 542462 75618 542546 75854
rect 542782 75618 578226 75854
rect 578462 75618 578546 75854
rect 578782 75618 585342 75854
rect 585578 75618 585662 75854
rect 585898 75618 592650 75854
rect -8726 75534 592650 75618
rect -8726 75298 -1974 75534
rect -1738 75298 -1654 75534
rect -1418 75298 2226 75534
rect 2462 75298 2546 75534
rect 2782 75298 38226 75534
rect 38462 75298 38546 75534
rect 38782 75298 74226 75534
rect 74462 75298 74546 75534
rect 74782 75298 110226 75534
rect 110462 75298 110546 75534
rect 110782 75298 146226 75534
rect 146462 75298 146546 75534
rect 146782 75298 182226 75534
rect 182462 75298 182546 75534
rect 182782 75298 218226 75534
rect 218462 75298 218546 75534
rect 218782 75298 254226 75534
rect 254462 75298 254546 75534
rect 254782 75298 290226 75534
rect 290462 75298 290546 75534
rect 290782 75298 326226 75534
rect 326462 75298 326546 75534
rect 326782 75298 362226 75534
rect 362462 75298 362546 75534
rect 362782 75298 398226 75534
rect 398462 75298 398546 75534
rect 398782 75298 434226 75534
rect 434462 75298 434546 75534
rect 434782 75298 470226 75534
rect 470462 75298 470546 75534
rect 470782 75298 506226 75534
rect 506462 75298 506546 75534
rect 506782 75298 542226 75534
rect 542462 75298 542546 75534
rect 542782 75298 578226 75534
rect 578462 75298 578546 75534
rect 578782 75298 585342 75534
rect 585578 75298 585662 75534
rect 585898 75298 592650 75534
rect -8726 75266 592650 75298
rect -8726 65894 592650 65926
rect -8726 65658 -8694 65894
rect -8458 65658 -8374 65894
rect -8138 65658 28266 65894
rect 28502 65658 28586 65894
rect 28822 65658 64266 65894
rect 64502 65658 64586 65894
rect 64822 65658 100266 65894
rect 100502 65658 100586 65894
rect 100822 65658 136266 65894
rect 136502 65658 136586 65894
rect 136822 65658 172266 65894
rect 172502 65658 172586 65894
rect 172822 65658 208266 65894
rect 208502 65658 208586 65894
rect 208822 65658 244266 65894
rect 244502 65658 244586 65894
rect 244822 65658 280266 65894
rect 280502 65658 280586 65894
rect 280822 65658 316266 65894
rect 316502 65658 316586 65894
rect 316822 65658 352266 65894
rect 352502 65658 352586 65894
rect 352822 65658 388266 65894
rect 388502 65658 388586 65894
rect 388822 65658 424266 65894
rect 424502 65658 424586 65894
rect 424822 65658 460266 65894
rect 460502 65658 460586 65894
rect 460822 65658 496266 65894
rect 496502 65658 496586 65894
rect 496822 65658 532266 65894
rect 532502 65658 532586 65894
rect 532822 65658 568266 65894
rect 568502 65658 568586 65894
rect 568822 65658 592062 65894
rect 592298 65658 592382 65894
rect 592618 65658 592650 65894
rect -8726 65574 592650 65658
rect -8726 65338 -8694 65574
rect -8458 65338 -8374 65574
rect -8138 65338 28266 65574
rect 28502 65338 28586 65574
rect 28822 65338 64266 65574
rect 64502 65338 64586 65574
rect 64822 65338 100266 65574
rect 100502 65338 100586 65574
rect 100822 65338 136266 65574
rect 136502 65338 136586 65574
rect 136822 65338 172266 65574
rect 172502 65338 172586 65574
rect 172822 65338 208266 65574
rect 208502 65338 208586 65574
rect 208822 65338 244266 65574
rect 244502 65338 244586 65574
rect 244822 65338 280266 65574
rect 280502 65338 280586 65574
rect 280822 65338 316266 65574
rect 316502 65338 316586 65574
rect 316822 65338 352266 65574
rect 352502 65338 352586 65574
rect 352822 65338 388266 65574
rect 388502 65338 388586 65574
rect 388822 65338 424266 65574
rect 424502 65338 424586 65574
rect 424822 65338 460266 65574
rect 460502 65338 460586 65574
rect 460822 65338 496266 65574
rect 496502 65338 496586 65574
rect 496822 65338 532266 65574
rect 532502 65338 532586 65574
rect 532822 65338 568266 65574
rect 568502 65338 568586 65574
rect 568822 65338 592062 65574
rect 592298 65338 592382 65574
rect 592618 65338 592650 65574
rect -8726 65306 592650 65338
rect -8726 62174 592650 62206
rect -8726 61938 -7734 62174
rect -7498 61938 -7414 62174
rect -7178 61938 24546 62174
rect 24782 61938 24866 62174
rect 25102 61938 60546 62174
rect 60782 61938 60866 62174
rect 61102 61938 96546 62174
rect 96782 61938 96866 62174
rect 97102 61938 132546 62174
rect 132782 61938 132866 62174
rect 133102 61938 168546 62174
rect 168782 61938 168866 62174
rect 169102 61938 204546 62174
rect 204782 61938 204866 62174
rect 205102 61938 240546 62174
rect 240782 61938 240866 62174
rect 241102 61938 276546 62174
rect 276782 61938 276866 62174
rect 277102 61938 312546 62174
rect 312782 61938 312866 62174
rect 313102 61938 348546 62174
rect 348782 61938 348866 62174
rect 349102 61938 384546 62174
rect 384782 61938 384866 62174
rect 385102 61938 420546 62174
rect 420782 61938 420866 62174
rect 421102 61938 456546 62174
rect 456782 61938 456866 62174
rect 457102 61938 492546 62174
rect 492782 61938 492866 62174
rect 493102 61938 528546 62174
rect 528782 61938 528866 62174
rect 529102 61938 564546 62174
rect 564782 61938 564866 62174
rect 565102 61938 591102 62174
rect 591338 61938 591422 62174
rect 591658 61938 592650 62174
rect -8726 61854 592650 61938
rect -8726 61618 -7734 61854
rect -7498 61618 -7414 61854
rect -7178 61618 24546 61854
rect 24782 61618 24866 61854
rect 25102 61618 60546 61854
rect 60782 61618 60866 61854
rect 61102 61618 96546 61854
rect 96782 61618 96866 61854
rect 97102 61618 132546 61854
rect 132782 61618 132866 61854
rect 133102 61618 168546 61854
rect 168782 61618 168866 61854
rect 169102 61618 204546 61854
rect 204782 61618 204866 61854
rect 205102 61618 240546 61854
rect 240782 61618 240866 61854
rect 241102 61618 276546 61854
rect 276782 61618 276866 61854
rect 277102 61618 312546 61854
rect 312782 61618 312866 61854
rect 313102 61618 348546 61854
rect 348782 61618 348866 61854
rect 349102 61618 384546 61854
rect 384782 61618 384866 61854
rect 385102 61618 420546 61854
rect 420782 61618 420866 61854
rect 421102 61618 456546 61854
rect 456782 61618 456866 61854
rect 457102 61618 492546 61854
rect 492782 61618 492866 61854
rect 493102 61618 528546 61854
rect 528782 61618 528866 61854
rect 529102 61618 564546 61854
rect 564782 61618 564866 61854
rect 565102 61618 591102 61854
rect 591338 61618 591422 61854
rect 591658 61618 592650 61854
rect -8726 61586 592650 61618
rect -8726 58454 592650 58486
rect -8726 58218 -6774 58454
rect -6538 58218 -6454 58454
rect -6218 58218 20826 58454
rect 21062 58218 21146 58454
rect 21382 58218 56826 58454
rect 57062 58218 57146 58454
rect 57382 58218 92826 58454
rect 93062 58218 93146 58454
rect 93382 58218 128826 58454
rect 129062 58218 129146 58454
rect 129382 58218 164826 58454
rect 165062 58218 165146 58454
rect 165382 58218 200826 58454
rect 201062 58218 201146 58454
rect 201382 58218 236826 58454
rect 237062 58218 237146 58454
rect 237382 58218 272826 58454
rect 273062 58218 273146 58454
rect 273382 58218 308826 58454
rect 309062 58218 309146 58454
rect 309382 58218 344826 58454
rect 345062 58218 345146 58454
rect 345382 58218 380826 58454
rect 381062 58218 381146 58454
rect 381382 58218 416826 58454
rect 417062 58218 417146 58454
rect 417382 58218 452826 58454
rect 453062 58218 453146 58454
rect 453382 58218 488826 58454
rect 489062 58218 489146 58454
rect 489382 58218 524826 58454
rect 525062 58218 525146 58454
rect 525382 58218 560826 58454
rect 561062 58218 561146 58454
rect 561382 58218 590142 58454
rect 590378 58218 590462 58454
rect 590698 58218 592650 58454
rect -8726 58134 592650 58218
rect -8726 57898 -6774 58134
rect -6538 57898 -6454 58134
rect -6218 57898 20826 58134
rect 21062 57898 21146 58134
rect 21382 57898 56826 58134
rect 57062 57898 57146 58134
rect 57382 57898 92826 58134
rect 93062 57898 93146 58134
rect 93382 57898 128826 58134
rect 129062 57898 129146 58134
rect 129382 57898 164826 58134
rect 165062 57898 165146 58134
rect 165382 57898 200826 58134
rect 201062 57898 201146 58134
rect 201382 57898 236826 58134
rect 237062 57898 237146 58134
rect 237382 57898 272826 58134
rect 273062 57898 273146 58134
rect 273382 57898 308826 58134
rect 309062 57898 309146 58134
rect 309382 57898 344826 58134
rect 345062 57898 345146 58134
rect 345382 57898 380826 58134
rect 381062 57898 381146 58134
rect 381382 57898 416826 58134
rect 417062 57898 417146 58134
rect 417382 57898 452826 58134
rect 453062 57898 453146 58134
rect 453382 57898 488826 58134
rect 489062 57898 489146 58134
rect 489382 57898 524826 58134
rect 525062 57898 525146 58134
rect 525382 57898 560826 58134
rect 561062 57898 561146 58134
rect 561382 57898 590142 58134
rect 590378 57898 590462 58134
rect 590698 57898 592650 58134
rect -8726 57866 592650 57898
rect -8726 54734 592650 54766
rect -8726 54498 -5814 54734
rect -5578 54498 -5494 54734
rect -5258 54498 17106 54734
rect 17342 54498 17426 54734
rect 17662 54498 53106 54734
rect 53342 54498 53426 54734
rect 53662 54498 89106 54734
rect 89342 54498 89426 54734
rect 89662 54498 125106 54734
rect 125342 54498 125426 54734
rect 125662 54498 161106 54734
rect 161342 54498 161426 54734
rect 161662 54498 197106 54734
rect 197342 54498 197426 54734
rect 197662 54498 233106 54734
rect 233342 54498 233426 54734
rect 233662 54498 269106 54734
rect 269342 54498 269426 54734
rect 269662 54498 305106 54734
rect 305342 54498 305426 54734
rect 305662 54498 341106 54734
rect 341342 54498 341426 54734
rect 341662 54498 377106 54734
rect 377342 54498 377426 54734
rect 377662 54498 413106 54734
rect 413342 54498 413426 54734
rect 413662 54498 449106 54734
rect 449342 54498 449426 54734
rect 449662 54498 485106 54734
rect 485342 54498 485426 54734
rect 485662 54498 521106 54734
rect 521342 54498 521426 54734
rect 521662 54498 557106 54734
rect 557342 54498 557426 54734
rect 557662 54498 589182 54734
rect 589418 54498 589502 54734
rect 589738 54498 592650 54734
rect -8726 54414 592650 54498
rect -8726 54178 -5814 54414
rect -5578 54178 -5494 54414
rect -5258 54178 17106 54414
rect 17342 54178 17426 54414
rect 17662 54178 53106 54414
rect 53342 54178 53426 54414
rect 53662 54178 89106 54414
rect 89342 54178 89426 54414
rect 89662 54178 125106 54414
rect 125342 54178 125426 54414
rect 125662 54178 161106 54414
rect 161342 54178 161426 54414
rect 161662 54178 197106 54414
rect 197342 54178 197426 54414
rect 197662 54178 233106 54414
rect 233342 54178 233426 54414
rect 233662 54178 269106 54414
rect 269342 54178 269426 54414
rect 269662 54178 305106 54414
rect 305342 54178 305426 54414
rect 305662 54178 341106 54414
rect 341342 54178 341426 54414
rect 341662 54178 377106 54414
rect 377342 54178 377426 54414
rect 377662 54178 413106 54414
rect 413342 54178 413426 54414
rect 413662 54178 449106 54414
rect 449342 54178 449426 54414
rect 449662 54178 485106 54414
rect 485342 54178 485426 54414
rect 485662 54178 521106 54414
rect 521342 54178 521426 54414
rect 521662 54178 557106 54414
rect 557342 54178 557426 54414
rect 557662 54178 589182 54414
rect 589418 54178 589502 54414
rect 589738 54178 592650 54414
rect -8726 54146 592650 54178
rect -8726 51014 592650 51046
rect -8726 50778 -4854 51014
rect -4618 50778 -4534 51014
rect -4298 50778 13386 51014
rect 13622 50778 13706 51014
rect 13942 50778 49386 51014
rect 49622 50778 49706 51014
rect 49942 50778 85386 51014
rect 85622 50778 85706 51014
rect 85942 50778 121386 51014
rect 121622 50778 121706 51014
rect 121942 50778 157386 51014
rect 157622 50778 157706 51014
rect 157942 50778 193386 51014
rect 193622 50778 193706 51014
rect 193942 50778 229386 51014
rect 229622 50778 229706 51014
rect 229942 50778 265386 51014
rect 265622 50778 265706 51014
rect 265942 50778 301386 51014
rect 301622 50778 301706 51014
rect 301942 50778 337386 51014
rect 337622 50778 337706 51014
rect 337942 50778 373386 51014
rect 373622 50778 373706 51014
rect 373942 50778 409386 51014
rect 409622 50778 409706 51014
rect 409942 50778 445386 51014
rect 445622 50778 445706 51014
rect 445942 50778 481386 51014
rect 481622 50778 481706 51014
rect 481942 50778 517386 51014
rect 517622 50778 517706 51014
rect 517942 50778 553386 51014
rect 553622 50778 553706 51014
rect 553942 50778 588222 51014
rect 588458 50778 588542 51014
rect 588778 50778 592650 51014
rect -8726 50694 592650 50778
rect -8726 50458 -4854 50694
rect -4618 50458 -4534 50694
rect -4298 50458 13386 50694
rect 13622 50458 13706 50694
rect 13942 50458 49386 50694
rect 49622 50458 49706 50694
rect 49942 50458 85386 50694
rect 85622 50458 85706 50694
rect 85942 50458 121386 50694
rect 121622 50458 121706 50694
rect 121942 50458 157386 50694
rect 157622 50458 157706 50694
rect 157942 50458 193386 50694
rect 193622 50458 193706 50694
rect 193942 50458 229386 50694
rect 229622 50458 229706 50694
rect 229942 50458 265386 50694
rect 265622 50458 265706 50694
rect 265942 50458 301386 50694
rect 301622 50458 301706 50694
rect 301942 50458 337386 50694
rect 337622 50458 337706 50694
rect 337942 50458 373386 50694
rect 373622 50458 373706 50694
rect 373942 50458 409386 50694
rect 409622 50458 409706 50694
rect 409942 50458 445386 50694
rect 445622 50458 445706 50694
rect 445942 50458 481386 50694
rect 481622 50458 481706 50694
rect 481942 50458 517386 50694
rect 517622 50458 517706 50694
rect 517942 50458 553386 50694
rect 553622 50458 553706 50694
rect 553942 50458 588222 50694
rect 588458 50458 588542 50694
rect 588778 50458 592650 50694
rect -8726 50426 592650 50458
rect -8726 47294 592650 47326
rect -8726 47058 -3894 47294
rect -3658 47058 -3574 47294
rect -3338 47058 9666 47294
rect 9902 47058 9986 47294
rect 10222 47058 45666 47294
rect 45902 47058 45986 47294
rect 46222 47058 81666 47294
rect 81902 47058 81986 47294
rect 82222 47058 117666 47294
rect 117902 47058 117986 47294
rect 118222 47058 153666 47294
rect 153902 47058 153986 47294
rect 154222 47058 189666 47294
rect 189902 47058 189986 47294
rect 190222 47058 225666 47294
rect 225902 47058 225986 47294
rect 226222 47058 261666 47294
rect 261902 47058 261986 47294
rect 262222 47058 297666 47294
rect 297902 47058 297986 47294
rect 298222 47058 333666 47294
rect 333902 47058 333986 47294
rect 334222 47058 369666 47294
rect 369902 47058 369986 47294
rect 370222 47058 405666 47294
rect 405902 47058 405986 47294
rect 406222 47058 441666 47294
rect 441902 47058 441986 47294
rect 442222 47058 477666 47294
rect 477902 47058 477986 47294
rect 478222 47058 513666 47294
rect 513902 47058 513986 47294
rect 514222 47058 549666 47294
rect 549902 47058 549986 47294
rect 550222 47058 587262 47294
rect 587498 47058 587582 47294
rect 587818 47058 592650 47294
rect -8726 46974 592650 47058
rect -8726 46738 -3894 46974
rect -3658 46738 -3574 46974
rect -3338 46738 9666 46974
rect 9902 46738 9986 46974
rect 10222 46738 45666 46974
rect 45902 46738 45986 46974
rect 46222 46738 81666 46974
rect 81902 46738 81986 46974
rect 82222 46738 117666 46974
rect 117902 46738 117986 46974
rect 118222 46738 153666 46974
rect 153902 46738 153986 46974
rect 154222 46738 189666 46974
rect 189902 46738 189986 46974
rect 190222 46738 225666 46974
rect 225902 46738 225986 46974
rect 226222 46738 261666 46974
rect 261902 46738 261986 46974
rect 262222 46738 297666 46974
rect 297902 46738 297986 46974
rect 298222 46738 333666 46974
rect 333902 46738 333986 46974
rect 334222 46738 369666 46974
rect 369902 46738 369986 46974
rect 370222 46738 405666 46974
rect 405902 46738 405986 46974
rect 406222 46738 441666 46974
rect 441902 46738 441986 46974
rect 442222 46738 477666 46974
rect 477902 46738 477986 46974
rect 478222 46738 513666 46974
rect 513902 46738 513986 46974
rect 514222 46738 549666 46974
rect 549902 46738 549986 46974
rect 550222 46738 587262 46974
rect 587498 46738 587582 46974
rect 587818 46738 592650 46974
rect -8726 46706 592650 46738
rect -8726 43574 592650 43606
rect -8726 43338 -2934 43574
rect -2698 43338 -2614 43574
rect -2378 43338 5946 43574
rect 6182 43338 6266 43574
rect 6502 43338 41946 43574
rect 42182 43338 42266 43574
rect 42502 43338 77946 43574
rect 78182 43338 78266 43574
rect 78502 43338 113946 43574
rect 114182 43338 114266 43574
rect 114502 43338 149946 43574
rect 150182 43338 150266 43574
rect 150502 43338 185946 43574
rect 186182 43338 186266 43574
rect 186502 43338 221946 43574
rect 222182 43338 222266 43574
rect 222502 43338 257946 43574
rect 258182 43338 258266 43574
rect 258502 43338 293946 43574
rect 294182 43338 294266 43574
rect 294502 43338 329946 43574
rect 330182 43338 330266 43574
rect 330502 43338 365946 43574
rect 366182 43338 366266 43574
rect 366502 43338 401946 43574
rect 402182 43338 402266 43574
rect 402502 43338 437946 43574
rect 438182 43338 438266 43574
rect 438502 43338 473946 43574
rect 474182 43338 474266 43574
rect 474502 43338 509946 43574
rect 510182 43338 510266 43574
rect 510502 43338 545946 43574
rect 546182 43338 546266 43574
rect 546502 43338 581946 43574
rect 582182 43338 582266 43574
rect 582502 43338 586302 43574
rect 586538 43338 586622 43574
rect 586858 43338 592650 43574
rect -8726 43254 592650 43338
rect -8726 43018 -2934 43254
rect -2698 43018 -2614 43254
rect -2378 43018 5946 43254
rect 6182 43018 6266 43254
rect 6502 43018 41946 43254
rect 42182 43018 42266 43254
rect 42502 43018 77946 43254
rect 78182 43018 78266 43254
rect 78502 43018 113946 43254
rect 114182 43018 114266 43254
rect 114502 43018 149946 43254
rect 150182 43018 150266 43254
rect 150502 43018 185946 43254
rect 186182 43018 186266 43254
rect 186502 43018 221946 43254
rect 222182 43018 222266 43254
rect 222502 43018 257946 43254
rect 258182 43018 258266 43254
rect 258502 43018 293946 43254
rect 294182 43018 294266 43254
rect 294502 43018 329946 43254
rect 330182 43018 330266 43254
rect 330502 43018 365946 43254
rect 366182 43018 366266 43254
rect 366502 43018 401946 43254
rect 402182 43018 402266 43254
rect 402502 43018 437946 43254
rect 438182 43018 438266 43254
rect 438502 43018 473946 43254
rect 474182 43018 474266 43254
rect 474502 43018 509946 43254
rect 510182 43018 510266 43254
rect 510502 43018 545946 43254
rect 546182 43018 546266 43254
rect 546502 43018 581946 43254
rect 582182 43018 582266 43254
rect 582502 43018 586302 43254
rect 586538 43018 586622 43254
rect 586858 43018 592650 43254
rect -8726 42986 592650 43018
rect -8726 39854 592650 39886
rect -8726 39618 -1974 39854
rect -1738 39618 -1654 39854
rect -1418 39618 2226 39854
rect 2462 39618 2546 39854
rect 2782 39618 38226 39854
rect 38462 39618 38546 39854
rect 38782 39618 74226 39854
rect 74462 39618 74546 39854
rect 74782 39618 110226 39854
rect 110462 39618 110546 39854
rect 110782 39618 146226 39854
rect 146462 39618 146546 39854
rect 146782 39618 182226 39854
rect 182462 39618 182546 39854
rect 182782 39618 218226 39854
rect 218462 39618 218546 39854
rect 218782 39618 254226 39854
rect 254462 39618 254546 39854
rect 254782 39618 290226 39854
rect 290462 39618 290546 39854
rect 290782 39618 326226 39854
rect 326462 39618 326546 39854
rect 326782 39618 362226 39854
rect 362462 39618 362546 39854
rect 362782 39618 398226 39854
rect 398462 39618 398546 39854
rect 398782 39618 434226 39854
rect 434462 39618 434546 39854
rect 434782 39618 470226 39854
rect 470462 39618 470546 39854
rect 470782 39618 506226 39854
rect 506462 39618 506546 39854
rect 506782 39618 542226 39854
rect 542462 39618 542546 39854
rect 542782 39618 578226 39854
rect 578462 39618 578546 39854
rect 578782 39618 585342 39854
rect 585578 39618 585662 39854
rect 585898 39618 592650 39854
rect -8726 39534 592650 39618
rect -8726 39298 -1974 39534
rect -1738 39298 -1654 39534
rect -1418 39298 2226 39534
rect 2462 39298 2546 39534
rect 2782 39298 38226 39534
rect 38462 39298 38546 39534
rect 38782 39298 74226 39534
rect 74462 39298 74546 39534
rect 74782 39298 110226 39534
rect 110462 39298 110546 39534
rect 110782 39298 146226 39534
rect 146462 39298 146546 39534
rect 146782 39298 182226 39534
rect 182462 39298 182546 39534
rect 182782 39298 218226 39534
rect 218462 39298 218546 39534
rect 218782 39298 254226 39534
rect 254462 39298 254546 39534
rect 254782 39298 290226 39534
rect 290462 39298 290546 39534
rect 290782 39298 326226 39534
rect 326462 39298 326546 39534
rect 326782 39298 362226 39534
rect 362462 39298 362546 39534
rect 362782 39298 398226 39534
rect 398462 39298 398546 39534
rect 398782 39298 434226 39534
rect 434462 39298 434546 39534
rect 434782 39298 470226 39534
rect 470462 39298 470546 39534
rect 470782 39298 506226 39534
rect 506462 39298 506546 39534
rect 506782 39298 542226 39534
rect 542462 39298 542546 39534
rect 542782 39298 578226 39534
rect 578462 39298 578546 39534
rect 578782 39298 585342 39534
rect 585578 39298 585662 39534
rect 585898 39298 592650 39534
rect -8726 39266 592650 39298
rect -8726 29894 592650 29926
rect -8726 29658 -8694 29894
rect -8458 29658 -8374 29894
rect -8138 29658 28266 29894
rect 28502 29658 28586 29894
rect 28822 29658 64266 29894
rect 64502 29658 64586 29894
rect 64822 29658 100266 29894
rect 100502 29658 100586 29894
rect 100822 29658 136266 29894
rect 136502 29658 136586 29894
rect 136822 29658 172266 29894
rect 172502 29658 172586 29894
rect 172822 29658 208266 29894
rect 208502 29658 208586 29894
rect 208822 29658 244266 29894
rect 244502 29658 244586 29894
rect 244822 29658 280266 29894
rect 280502 29658 280586 29894
rect 280822 29658 316266 29894
rect 316502 29658 316586 29894
rect 316822 29658 352266 29894
rect 352502 29658 352586 29894
rect 352822 29658 388266 29894
rect 388502 29658 388586 29894
rect 388822 29658 424266 29894
rect 424502 29658 424586 29894
rect 424822 29658 460266 29894
rect 460502 29658 460586 29894
rect 460822 29658 496266 29894
rect 496502 29658 496586 29894
rect 496822 29658 532266 29894
rect 532502 29658 532586 29894
rect 532822 29658 568266 29894
rect 568502 29658 568586 29894
rect 568822 29658 592062 29894
rect 592298 29658 592382 29894
rect 592618 29658 592650 29894
rect -8726 29574 592650 29658
rect -8726 29338 -8694 29574
rect -8458 29338 -8374 29574
rect -8138 29338 28266 29574
rect 28502 29338 28586 29574
rect 28822 29338 64266 29574
rect 64502 29338 64586 29574
rect 64822 29338 100266 29574
rect 100502 29338 100586 29574
rect 100822 29338 136266 29574
rect 136502 29338 136586 29574
rect 136822 29338 172266 29574
rect 172502 29338 172586 29574
rect 172822 29338 208266 29574
rect 208502 29338 208586 29574
rect 208822 29338 244266 29574
rect 244502 29338 244586 29574
rect 244822 29338 280266 29574
rect 280502 29338 280586 29574
rect 280822 29338 316266 29574
rect 316502 29338 316586 29574
rect 316822 29338 352266 29574
rect 352502 29338 352586 29574
rect 352822 29338 388266 29574
rect 388502 29338 388586 29574
rect 388822 29338 424266 29574
rect 424502 29338 424586 29574
rect 424822 29338 460266 29574
rect 460502 29338 460586 29574
rect 460822 29338 496266 29574
rect 496502 29338 496586 29574
rect 496822 29338 532266 29574
rect 532502 29338 532586 29574
rect 532822 29338 568266 29574
rect 568502 29338 568586 29574
rect 568822 29338 592062 29574
rect 592298 29338 592382 29574
rect 592618 29338 592650 29574
rect -8726 29306 592650 29338
rect -8726 26174 592650 26206
rect -8726 25938 -7734 26174
rect -7498 25938 -7414 26174
rect -7178 25938 24546 26174
rect 24782 25938 24866 26174
rect 25102 25938 60546 26174
rect 60782 25938 60866 26174
rect 61102 25938 96546 26174
rect 96782 25938 96866 26174
rect 97102 25938 132546 26174
rect 132782 25938 132866 26174
rect 133102 25938 168546 26174
rect 168782 25938 168866 26174
rect 169102 25938 204546 26174
rect 204782 25938 204866 26174
rect 205102 25938 240546 26174
rect 240782 25938 240866 26174
rect 241102 25938 276546 26174
rect 276782 25938 276866 26174
rect 277102 25938 312546 26174
rect 312782 25938 312866 26174
rect 313102 25938 348546 26174
rect 348782 25938 348866 26174
rect 349102 25938 384546 26174
rect 384782 25938 384866 26174
rect 385102 25938 420546 26174
rect 420782 25938 420866 26174
rect 421102 25938 456546 26174
rect 456782 25938 456866 26174
rect 457102 25938 492546 26174
rect 492782 25938 492866 26174
rect 493102 25938 528546 26174
rect 528782 25938 528866 26174
rect 529102 25938 564546 26174
rect 564782 25938 564866 26174
rect 565102 25938 591102 26174
rect 591338 25938 591422 26174
rect 591658 25938 592650 26174
rect -8726 25854 592650 25938
rect -8726 25618 -7734 25854
rect -7498 25618 -7414 25854
rect -7178 25618 24546 25854
rect 24782 25618 24866 25854
rect 25102 25618 60546 25854
rect 60782 25618 60866 25854
rect 61102 25618 96546 25854
rect 96782 25618 96866 25854
rect 97102 25618 132546 25854
rect 132782 25618 132866 25854
rect 133102 25618 168546 25854
rect 168782 25618 168866 25854
rect 169102 25618 204546 25854
rect 204782 25618 204866 25854
rect 205102 25618 240546 25854
rect 240782 25618 240866 25854
rect 241102 25618 276546 25854
rect 276782 25618 276866 25854
rect 277102 25618 312546 25854
rect 312782 25618 312866 25854
rect 313102 25618 348546 25854
rect 348782 25618 348866 25854
rect 349102 25618 384546 25854
rect 384782 25618 384866 25854
rect 385102 25618 420546 25854
rect 420782 25618 420866 25854
rect 421102 25618 456546 25854
rect 456782 25618 456866 25854
rect 457102 25618 492546 25854
rect 492782 25618 492866 25854
rect 493102 25618 528546 25854
rect 528782 25618 528866 25854
rect 529102 25618 564546 25854
rect 564782 25618 564866 25854
rect 565102 25618 591102 25854
rect 591338 25618 591422 25854
rect 591658 25618 592650 25854
rect -8726 25586 592650 25618
rect -8726 22454 592650 22486
rect -8726 22218 -6774 22454
rect -6538 22218 -6454 22454
rect -6218 22218 20826 22454
rect 21062 22218 21146 22454
rect 21382 22218 56826 22454
rect 57062 22218 57146 22454
rect 57382 22218 92826 22454
rect 93062 22218 93146 22454
rect 93382 22218 128826 22454
rect 129062 22218 129146 22454
rect 129382 22218 164826 22454
rect 165062 22218 165146 22454
rect 165382 22218 200826 22454
rect 201062 22218 201146 22454
rect 201382 22218 236826 22454
rect 237062 22218 237146 22454
rect 237382 22218 272826 22454
rect 273062 22218 273146 22454
rect 273382 22218 308826 22454
rect 309062 22218 309146 22454
rect 309382 22218 344826 22454
rect 345062 22218 345146 22454
rect 345382 22218 380826 22454
rect 381062 22218 381146 22454
rect 381382 22218 416826 22454
rect 417062 22218 417146 22454
rect 417382 22218 452826 22454
rect 453062 22218 453146 22454
rect 453382 22218 488826 22454
rect 489062 22218 489146 22454
rect 489382 22218 524826 22454
rect 525062 22218 525146 22454
rect 525382 22218 560826 22454
rect 561062 22218 561146 22454
rect 561382 22218 590142 22454
rect 590378 22218 590462 22454
rect 590698 22218 592650 22454
rect -8726 22134 592650 22218
rect -8726 21898 -6774 22134
rect -6538 21898 -6454 22134
rect -6218 21898 20826 22134
rect 21062 21898 21146 22134
rect 21382 21898 56826 22134
rect 57062 21898 57146 22134
rect 57382 21898 92826 22134
rect 93062 21898 93146 22134
rect 93382 21898 128826 22134
rect 129062 21898 129146 22134
rect 129382 21898 164826 22134
rect 165062 21898 165146 22134
rect 165382 21898 200826 22134
rect 201062 21898 201146 22134
rect 201382 21898 236826 22134
rect 237062 21898 237146 22134
rect 237382 21898 272826 22134
rect 273062 21898 273146 22134
rect 273382 21898 308826 22134
rect 309062 21898 309146 22134
rect 309382 21898 344826 22134
rect 345062 21898 345146 22134
rect 345382 21898 380826 22134
rect 381062 21898 381146 22134
rect 381382 21898 416826 22134
rect 417062 21898 417146 22134
rect 417382 21898 452826 22134
rect 453062 21898 453146 22134
rect 453382 21898 488826 22134
rect 489062 21898 489146 22134
rect 489382 21898 524826 22134
rect 525062 21898 525146 22134
rect 525382 21898 560826 22134
rect 561062 21898 561146 22134
rect 561382 21898 590142 22134
rect 590378 21898 590462 22134
rect 590698 21898 592650 22134
rect -8726 21866 592650 21898
rect -8726 18734 592650 18766
rect -8726 18498 -5814 18734
rect -5578 18498 -5494 18734
rect -5258 18498 17106 18734
rect 17342 18498 17426 18734
rect 17662 18498 53106 18734
rect 53342 18498 53426 18734
rect 53662 18498 89106 18734
rect 89342 18498 89426 18734
rect 89662 18498 125106 18734
rect 125342 18498 125426 18734
rect 125662 18498 161106 18734
rect 161342 18498 161426 18734
rect 161662 18498 197106 18734
rect 197342 18498 197426 18734
rect 197662 18498 233106 18734
rect 233342 18498 233426 18734
rect 233662 18498 269106 18734
rect 269342 18498 269426 18734
rect 269662 18498 305106 18734
rect 305342 18498 305426 18734
rect 305662 18498 341106 18734
rect 341342 18498 341426 18734
rect 341662 18498 377106 18734
rect 377342 18498 377426 18734
rect 377662 18498 413106 18734
rect 413342 18498 413426 18734
rect 413662 18498 449106 18734
rect 449342 18498 449426 18734
rect 449662 18498 485106 18734
rect 485342 18498 485426 18734
rect 485662 18498 521106 18734
rect 521342 18498 521426 18734
rect 521662 18498 557106 18734
rect 557342 18498 557426 18734
rect 557662 18498 589182 18734
rect 589418 18498 589502 18734
rect 589738 18498 592650 18734
rect -8726 18414 592650 18498
rect -8726 18178 -5814 18414
rect -5578 18178 -5494 18414
rect -5258 18178 17106 18414
rect 17342 18178 17426 18414
rect 17662 18178 53106 18414
rect 53342 18178 53426 18414
rect 53662 18178 89106 18414
rect 89342 18178 89426 18414
rect 89662 18178 125106 18414
rect 125342 18178 125426 18414
rect 125662 18178 161106 18414
rect 161342 18178 161426 18414
rect 161662 18178 197106 18414
rect 197342 18178 197426 18414
rect 197662 18178 233106 18414
rect 233342 18178 233426 18414
rect 233662 18178 269106 18414
rect 269342 18178 269426 18414
rect 269662 18178 305106 18414
rect 305342 18178 305426 18414
rect 305662 18178 341106 18414
rect 341342 18178 341426 18414
rect 341662 18178 377106 18414
rect 377342 18178 377426 18414
rect 377662 18178 413106 18414
rect 413342 18178 413426 18414
rect 413662 18178 449106 18414
rect 449342 18178 449426 18414
rect 449662 18178 485106 18414
rect 485342 18178 485426 18414
rect 485662 18178 521106 18414
rect 521342 18178 521426 18414
rect 521662 18178 557106 18414
rect 557342 18178 557426 18414
rect 557662 18178 589182 18414
rect 589418 18178 589502 18414
rect 589738 18178 592650 18414
rect -8726 18146 592650 18178
rect -8726 15014 592650 15046
rect -8726 14778 -4854 15014
rect -4618 14778 -4534 15014
rect -4298 14778 13386 15014
rect 13622 14778 13706 15014
rect 13942 14778 49386 15014
rect 49622 14778 49706 15014
rect 49942 14778 85386 15014
rect 85622 14778 85706 15014
rect 85942 14778 121386 15014
rect 121622 14778 121706 15014
rect 121942 14778 157386 15014
rect 157622 14778 157706 15014
rect 157942 14778 193386 15014
rect 193622 14778 193706 15014
rect 193942 14778 229386 15014
rect 229622 14778 229706 15014
rect 229942 14778 265386 15014
rect 265622 14778 265706 15014
rect 265942 14778 301386 15014
rect 301622 14778 301706 15014
rect 301942 14778 337386 15014
rect 337622 14778 337706 15014
rect 337942 14778 373386 15014
rect 373622 14778 373706 15014
rect 373942 14778 409386 15014
rect 409622 14778 409706 15014
rect 409942 14778 445386 15014
rect 445622 14778 445706 15014
rect 445942 14778 481386 15014
rect 481622 14778 481706 15014
rect 481942 14778 517386 15014
rect 517622 14778 517706 15014
rect 517942 14778 553386 15014
rect 553622 14778 553706 15014
rect 553942 14778 588222 15014
rect 588458 14778 588542 15014
rect 588778 14778 592650 15014
rect -8726 14694 592650 14778
rect -8726 14458 -4854 14694
rect -4618 14458 -4534 14694
rect -4298 14458 13386 14694
rect 13622 14458 13706 14694
rect 13942 14458 49386 14694
rect 49622 14458 49706 14694
rect 49942 14458 85386 14694
rect 85622 14458 85706 14694
rect 85942 14458 121386 14694
rect 121622 14458 121706 14694
rect 121942 14458 157386 14694
rect 157622 14458 157706 14694
rect 157942 14458 193386 14694
rect 193622 14458 193706 14694
rect 193942 14458 229386 14694
rect 229622 14458 229706 14694
rect 229942 14458 265386 14694
rect 265622 14458 265706 14694
rect 265942 14458 301386 14694
rect 301622 14458 301706 14694
rect 301942 14458 337386 14694
rect 337622 14458 337706 14694
rect 337942 14458 373386 14694
rect 373622 14458 373706 14694
rect 373942 14458 409386 14694
rect 409622 14458 409706 14694
rect 409942 14458 445386 14694
rect 445622 14458 445706 14694
rect 445942 14458 481386 14694
rect 481622 14458 481706 14694
rect 481942 14458 517386 14694
rect 517622 14458 517706 14694
rect 517942 14458 553386 14694
rect 553622 14458 553706 14694
rect 553942 14458 588222 14694
rect 588458 14458 588542 14694
rect 588778 14458 592650 14694
rect -8726 14426 592650 14458
rect 57708 12018 191612 12060
rect 57708 11782 57750 12018
rect 57986 11782 191334 12018
rect 191570 11782 191612 12018
rect 57708 11740 191612 11782
rect -8726 11294 592650 11326
rect -8726 11058 -3894 11294
rect -3658 11058 -3574 11294
rect -3338 11058 9666 11294
rect 9902 11058 9986 11294
rect 10222 11058 45666 11294
rect 45902 11058 45986 11294
rect 46222 11058 81666 11294
rect 81902 11058 81986 11294
rect 82222 11058 117666 11294
rect 117902 11058 117986 11294
rect 118222 11058 153666 11294
rect 153902 11058 153986 11294
rect 154222 11058 189666 11294
rect 189902 11058 189986 11294
rect 190222 11058 225666 11294
rect 225902 11058 225986 11294
rect 226222 11058 261666 11294
rect 261902 11058 261986 11294
rect 262222 11058 297666 11294
rect 297902 11058 297986 11294
rect 298222 11058 333666 11294
rect 333902 11058 333986 11294
rect 334222 11058 369666 11294
rect 369902 11058 369986 11294
rect 370222 11058 405666 11294
rect 405902 11058 405986 11294
rect 406222 11058 441666 11294
rect 441902 11058 441986 11294
rect 442222 11058 477666 11294
rect 477902 11058 477986 11294
rect 478222 11058 513666 11294
rect 513902 11058 513986 11294
rect 514222 11058 549666 11294
rect 549902 11058 549986 11294
rect 550222 11058 587262 11294
rect 587498 11058 587582 11294
rect 587818 11058 592650 11294
rect -8726 10974 592650 11058
rect -8726 10738 -3894 10974
rect -3658 10738 -3574 10974
rect -3338 10738 9666 10974
rect 9902 10738 9986 10974
rect 10222 10738 45666 10974
rect 45902 10738 45986 10974
rect 46222 10738 81666 10974
rect 81902 10738 81986 10974
rect 82222 10738 117666 10974
rect 117902 10738 117986 10974
rect 118222 10738 153666 10974
rect 153902 10738 153986 10974
rect 154222 10738 189666 10974
rect 189902 10738 189986 10974
rect 190222 10738 225666 10974
rect 225902 10738 225986 10974
rect 226222 10738 261666 10974
rect 261902 10738 261986 10974
rect 262222 10738 297666 10974
rect 297902 10738 297986 10974
rect 298222 10738 333666 10974
rect 333902 10738 333986 10974
rect 334222 10738 369666 10974
rect 369902 10738 369986 10974
rect 370222 10738 405666 10974
rect 405902 10738 405986 10974
rect 406222 10738 441666 10974
rect 441902 10738 441986 10974
rect 442222 10738 477666 10974
rect 477902 10738 477986 10974
rect 478222 10738 513666 10974
rect 513902 10738 513986 10974
rect 514222 10738 549666 10974
rect 549902 10738 549986 10974
rect 550222 10738 587262 10974
rect 587498 10738 587582 10974
rect 587818 10738 592650 10974
rect -8726 10706 592650 10738
rect 27716 9978 145244 10020
rect 27716 9742 27758 9978
rect 27994 9742 144966 9978
rect 145202 9742 145244 9978
rect 27716 9700 145244 9742
rect 412460 9298 431916 9340
rect 412460 9062 431638 9298
rect 431874 9062 431916 9298
rect 412460 9020 431916 9062
rect 412460 8660 412780 9020
rect 67276 8618 163092 8660
rect 67276 8382 67318 8618
rect 67554 8382 162814 8618
rect 163050 8382 163092 8618
rect 67276 8340 163092 8382
rect 296540 8618 412780 8660
rect 296540 8382 296582 8618
rect 296818 8382 412780 8618
rect 296540 8340 412780 8382
rect -8726 7574 592650 7606
rect -8726 7338 -2934 7574
rect -2698 7338 -2614 7574
rect -2378 7338 5946 7574
rect 6182 7338 6266 7574
rect 6502 7338 41946 7574
rect 42182 7338 42266 7574
rect 42502 7338 77946 7574
rect 78182 7338 78266 7574
rect 78502 7338 113946 7574
rect 114182 7338 114266 7574
rect 114502 7338 149946 7574
rect 150182 7338 150266 7574
rect 150502 7338 185946 7574
rect 186182 7338 186266 7574
rect 186502 7338 221946 7574
rect 222182 7338 222266 7574
rect 222502 7338 257946 7574
rect 258182 7338 258266 7574
rect 258502 7338 293946 7574
rect 294182 7338 294266 7574
rect 294502 7338 329946 7574
rect 330182 7338 330266 7574
rect 330502 7338 365946 7574
rect 366182 7338 366266 7574
rect 366502 7338 401946 7574
rect 402182 7338 402266 7574
rect 402502 7338 437946 7574
rect 438182 7338 438266 7574
rect 438502 7338 473946 7574
rect 474182 7338 474266 7574
rect 474502 7338 509946 7574
rect 510182 7338 510266 7574
rect 510502 7338 545946 7574
rect 546182 7338 546266 7574
rect 546502 7338 581946 7574
rect 582182 7338 582266 7574
rect 582502 7338 586302 7574
rect 586538 7338 586622 7574
rect 586858 7338 592650 7574
rect -8726 7254 592650 7338
rect -8726 7018 -2934 7254
rect -2698 7018 -2614 7254
rect -2378 7018 5946 7254
rect 6182 7018 6266 7254
rect 6502 7018 41946 7254
rect 42182 7018 42266 7254
rect 42502 7018 77946 7254
rect 78182 7018 78266 7254
rect 78502 7018 113946 7254
rect 114182 7018 114266 7254
rect 114502 7018 149946 7254
rect 150182 7018 150266 7254
rect 150502 7018 185946 7254
rect 186182 7018 186266 7254
rect 186502 7018 221946 7254
rect 222182 7018 222266 7254
rect 222502 7018 257946 7254
rect 258182 7018 258266 7254
rect 258502 7018 293946 7254
rect 294182 7018 294266 7254
rect 294502 7018 329946 7254
rect 330182 7018 330266 7254
rect 330502 7018 365946 7254
rect 366182 7018 366266 7254
rect 366502 7018 401946 7254
rect 402182 7018 402266 7254
rect 402502 7018 437946 7254
rect 438182 7018 438266 7254
rect 438502 7018 473946 7254
rect 474182 7018 474266 7254
rect 474502 7018 509946 7254
rect 510182 7018 510266 7254
rect 510502 7018 545946 7254
rect 546182 7018 546266 7254
rect 546502 7018 581946 7254
rect 582182 7018 582266 7254
rect 582502 7018 586302 7254
rect 586538 7018 586622 7254
rect 586858 7018 592650 7254
rect -8726 6986 592650 7018
rect 191660 6578 339180 6620
rect 191660 6342 191702 6578
rect 191938 6342 338902 6578
rect 339138 6342 339180 6578
rect 191660 6300 339180 6342
rect 43908 5898 190876 5940
rect 43908 5662 43950 5898
rect 44186 5662 190598 5898
rect 190834 5662 190876 5898
rect 43908 5620 190876 5662
rect 180620 5218 191612 5260
rect 180620 4982 191334 5218
rect 191570 4982 191612 5218
rect 180620 4940 191612 4982
rect 180620 4580 180940 4940
rect 12260 4538 91332 4580
rect 12260 4302 12302 4538
rect 12538 4302 91054 4538
rect 91290 4302 91332 4538
rect 12260 4260 91332 4302
rect 113460 4538 180940 4580
rect 113460 4302 113502 4538
rect 113738 4302 180940 4538
rect 113460 4260 180940 4302
rect 203988 4538 338628 4580
rect 203988 4302 204030 4538
rect 204266 4302 338350 4538
rect 338586 4302 338628 4538
rect 203988 4260 338628 4302
rect -8726 3854 592650 3886
rect -8726 3618 -1974 3854
rect -1738 3618 -1654 3854
rect -1418 3618 2226 3854
rect 2462 3618 2546 3854
rect 2782 3618 38226 3854
rect 38462 3618 38546 3854
rect 38782 3618 74226 3854
rect 74462 3618 74546 3854
rect 74782 3618 110226 3854
rect 110462 3618 110546 3854
rect 110782 3618 146226 3854
rect 146462 3618 146546 3854
rect 146782 3618 182226 3854
rect 182462 3618 182546 3854
rect 182782 3618 218226 3854
rect 218462 3618 218546 3854
rect 218782 3618 254226 3854
rect 254462 3618 254546 3854
rect 254782 3618 290226 3854
rect 290462 3618 290546 3854
rect 290782 3618 326226 3854
rect 326462 3618 326546 3854
rect 326782 3618 362226 3854
rect 362462 3618 362546 3854
rect 362782 3618 398226 3854
rect 398462 3618 398546 3854
rect 398782 3618 434226 3854
rect 434462 3618 434546 3854
rect 434782 3618 470226 3854
rect 470462 3618 470546 3854
rect 470782 3618 506226 3854
rect 506462 3618 506546 3854
rect 506782 3618 542226 3854
rect 542462 3618 542546 3854
rect 542782 3618 578226 3854
rect 578462 3618 578546 3854
rect 578782 3618 585342 3854
rect 585578 3618 585662 3854
rect 585898 3618 592650 3854
rect -8726 3534 592650 3618
rect -8726 3298 -1974 3534
rect -1738 3298 -1654 3534
rect -1418 3298 2226 3534
rect 2462 3298 2546 3534
rect 2782 3298 38226 3534
rect 38462 3298 38546 3534
rect 38782 3298 74226 3534
rect 74462 3298 74546 3534
rect 74782 3298 110226 3534
rect 110462 3298 110546 3534
rect 110782 3298 146226 3534
rect 146462 3298 146546 3534
rect 146782 3298 182226 3534
rect 182462 3298 182546 3534
rect 182782 3298 218226 3534
rect 218462 3298 218546 3534
rect 218782 3298 254226 3534
rect 254462 3298 254546 3534
rect 254782 3298 290226 3534
rect 290462 3298 290546 3534
rect 290782 3298 326226 3534
rect 326462 3298 326546 3534
rect 326782 3298 362226 3534
rect 362462 3298 362546 3534
rect 362782 3298 398226 3534
rect 398462 3298 398546 3534
rect 398782 3298 434226 3534
rect 434462 3298 434546 3534
rect 434782 3298 470226 3534
rect 470462 3298 470546 3534
rect 470782 3298 506226 3534
rect 506462 3298 506546 3534
rect 506782 3298 542226 3534
rect 542462 3298 542546 3534
rect 542782 3298 578226 3534
rect 578462 3298 578546 3534
rect 578782 3298 585342 3534
rect 585578 3298 585662 3534
rect 585898 3298 592650 3534
rect -8726 3266 592650 3298
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 2226 -346
rect 2462 -582 2546 -346
rect 2782 -582 38226 -346
rect 38462 -582 38546 -346
rect 38782 -582 74226 -346
rect 74462 -582 74546 -346
rect 74782 -582 110226 -346
rect 110462 -582 110546 -346
rect 110782 -582 146226 -346
rect 146462 -582 146546 -346
rect 146782 -582 182226 -346
rect 182462 -582 182546 -346
rect 182782 -582 218226 -346
rect 218462 -582 218546 -346
rect 218782 -582 254226 -346
rect 254462 -582 254546 -346
rect 254782 -582 290226 -346
rect 290462 -582 290546 -346
rect 290782 -582 326226 -346
rect 326462 -582 326546 -346
rect 326782 -582 362226 -346
rect 362462 -582 362546 -346
rect 362782 -582 398226 -346
rect 398462 -582 398546 -346
rect 398782 -582 434226 -346
rect 434462 -582 434546 -346
rect 434782 -582 470226 -346
rect 470462 -582 470546 -346
rect 470782 -582 506226 -346
rect 506462 -582 506546 -346
rect 506782 -582 542226 -346
rect 542462 -582 542546 -346
rect 542782 -582 578226 -346
rect 578462 -582 578546 -346
rect 578782 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 2226 -666
rect 2462 -902 2546 -666
rect 2782 -902 38226 -666
rect 38462 -902 38546 -666
rect 38782 -902 74226 -666
rect 74462 -902 74546 -666
rect 74782 -902 110226 -666
rect 110462 -902 110546 -666
rect 110782 -902 146226 -666
rect 146462 -902 146546 -666
rect 146782 -902 182226 -666
rect 182462 -902 182546 -666
rect 182782 -902 218226 -666
rect 218462 -902 218546 -666
rect 218782 -902 254226 -666
rect 254462 -902 254546 -666
rect 254782 -902 290226 -666
rect 290462 -902 290546 -666
rect 290782 -902 326226 -666
rect 326462 -902 326546 -666
rect 326782 -902 362226 -666
rect 362462 -902 362546 -666
rect 362782 -902 398226 -666
rect 398462 -902 398546 -666
rect 398782 -902 434226 -666
rect 434462 -902 434546 -666
rect 434782 -902 470226 -666
rect 470462 -902 470546 -666
rect 470782 -902 506226 -666
rect 506462 -902 506546 -666
rect 506782 -902 542226 -666
rect 542462 -902 542546 -666
rect 542782 -902 578226 -666
rect 578462 -902 578546 -666
rect 578782 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5946 -1306
rect 6182 -1542 6266 -1306
rect 6502 -1542 41946 -1306
rect 42182 -1542 42266 -1306
rect 42502 -1542 77946 -1306
rect 78182 -1542 78266 -1306
rect 78502 -1542 113946 -1306
rect 114182 -1542 114266 -1306
rect 114502 -1542 149946 -1306
rect 150182 -1542 150266 -1306
rect 150502 -1542 185946 -1306
rect 186182 -1542 186266 -1306
rect 186502 -1542 221946 -1306
rect 222182 -1542 222266 -1306
rect 222502 -1542 257946 -1306
rect 258182 -1542 258266 -1306
rect 258502 -1542 293946 -1306
rect 294182 -1542 294266 -1306
rect 294502 -1542 329946 -1306
rect 330182 -1542 330266 -1306
rect 330502 -1542 365946 -1306
rect 366182 -1542 366266 -1306
rect 366502 -1542 401946 -1306
rect 402182 -1542 402266 -1306
rect 402502 -1542 437946 -1306
rect 438182 -1542 438266 -1306
rect 438502 -1542 473946 -1306
rect 474182 -1542 474266 -1306
rect 474502 -1542 509946 -1306
rect 510182 -1542 510266 -1306
rect 510502 -1542 545946 -1306
rect 546182 -1542 546266 -1306
rect 546502 -1542 581946 -1306
rect 582182 -1542 582266 -1306
rect 582502 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5946 -1626
rect 6182 -1862 6266 -1626
rect 6502 -1862 41946 -1626
rect 42182 -1862 42266 -1626
rect 42502 -1862 77946 -1626
rect 78182 -1862 78266 -1626
rect 78502 -1862 113946 -1626
rect 114182 -1862 114266 -1626
rect 114502 -1862 149946 -1626
rect 150182 -1862 150266 -1626
rect 150502 -1862 185946 -1626
rect 186182 -1862 186266 -1626
rect 186502 -1862 221946 -1626
rect 222182 -1862 222266 -1626
rect 222502 -1862 257946 -1626
rect 258182 -1862 258266 -1626
rect 258502 -1862 293946 -1626
rect 294182 -1862 294266 -1626
rect 294502 -1862 329946 -1626
rect 330182 -1862 330266 -1626
rect 330502 -1862 365946 -1626
rect 366182 -1862 366266 -1626
rect 366502 -1862 401946 -1626
rect 402182 -1862 402266 -1626
rect 402502 -1862 437946 -1626
rect 438182 -1862 438266 -1626
rect 438502 -1862 473946 -1626
rect 474182 -1862 474266 -1626
rect 474502 -1862 509946 -1626
rect 510182 -1862 510266 -1626
rect 510502 -1862 545946 -1626
rect 546182 -1862 546266 -1626
rect 546502 -1862 581946 -1626
rect 582182 -1862 582266 -1626
rect 582502 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9666 -2266
rect 9902 -2502 9986 -2266
rect 10222 -2502 45666 -2266
rect 45902 -2502 45986 -2266
rect 46222 -2502 81666 -2266
rect 81902 -2502 81986 -2266
rect 82222 -2502 117666 -2266
rect 117902 -2502 117986 -2266
rect 118222 -2502 153666 -2266
rect 153902 -2502 153986 -2266
rect 154222 -2502 189666 -2266
rect 189902 -2502 189986 -2266
rect 190222 -2502 225666 -2266
rect 225902 -2502 225986 -2266
rect 226222 -2502 261666 -2266
rect 261902 -2502 261986 -2266
rect 262222 -2502 297666 -2266
rect 297902 -2502 297986 -2266
rect 298222 -2502 333666 -2266
rect 333902 -2502 333986 -2266
rect 334222 -2502 369666 -2266
rect 369902 -2502 369986 -2266
rect 370222 -2502 405666 -2266
rect 405902 -2502 405986 -2266
rect 406222 -2502 441666 -2266
rect 441902 -2502 441986 -2266
rect 442222 -2502 477666 -2266
rect 477902 -2502 477986 -2266
rect 478222 -2502 513666 -2266
rect 513902 -2502 513986 -2266
rect 514222 -2502 549666 -2266
rect 549902 -2502 549986 -2266
rect 550222 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9666 -2586
rect 9902 -2822 9986 -2586
rect 10222 -2822 45666 -2586
rect 45902 -2822 45986 -2586
rect 46222 -2822 81666 -2586
rect 81902 -2822 81986 -2586
rect 82222 -2822 117666 -2586
rect 117902 -2822 117986 -2586
rect 118222 -2822 153666 -2586
rect 153902 -2822 153986 -2586
rect 154222 -2822 189666 -2586
rect 189902 -2822 189986 -2586
rect 190222 -2822 225666 -2586
rect 225902 -2822 225986 -2586
rect 226222 -2822 261666 -2586
rect 261902 -2822 261986 -2586
rect 262222 -2822 297666 -2586
rect 297902 -2822 297986 -2586
rect 298222 -2822 333666 -2586
rect 333902 -2822 333986 -2586
rect 334222 -2822 369666 -2586
rect 369902 -2822 369986 -2586
rect 370222 -2822 405666 -2586
rect 405902 -2822 405986 -2586
rect 406222 -2822 441666 -2586
rect 441902 -2822 441986 -2586
rect 442222 -2822 477666 -2586
rect 477902 -2822 477986 -2586
rect 478222 -2822 513666 -2586
rect 513902 -2822 513986 -2586
rect 514222 -2822 549666 -2586
rect 549902 -2822 549986 -2586
rect 550222 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 13386 -3226
rect 13622 -3462 13706 -3226
rect 13942 -3462 49386 -3226
rect 49622 -3462 49706 -3226
rect 49942 -3462 85386 -3226
rect 85622 -3462 85706 -3226
rect 85942 -3462 121386 -3226
rect 121622 -3462 121706 -3226
rect 121942 -3462 157386 -3226
rect 157622 -3462 157706 -3226
rect 157942 -3462 193386 -3226
rect 193622 -3462 193706 -3226
rect 193942 -3462 229386 -3226
rect 229622 -3462 229706 -3226
rect 229942 -3462 265386 -3226
rect 265622 -3462 265706 -3226
rect 265942 -3462 301386 -3226
rect 301622 -3462 301706 -3226
rect 301942 -3462 337386 -3226
rect 337622 -3462 337706 -3226
rect 337942 -3462 373386 -3226
rect 373622 -3462 373706 -3226
rect 373942 -3462 409386 -3226
rect 409622 -3462 409706 -3226
rect 409942 -3462 445386 -3226
rect 445622 -3462 445706 -3226
rect 445942 -3462 481386 -3226
rect 481622 -3462 481706 -3226
rect 481942 -3462 517386 -3226
rect 517622 -3462 517706 -3226
rect 517942 -3462 553386 -3226
rect 553622 -3462 553706 -3226
rect 553942 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 13386 -3546
rect 13622 -3782 13706 -3546
rect 13942 -3782 49386 -3546
rect 49622 -3782 49706 -3546
rect 49942 -3782 85386 -3546
rect 85622 -3782 85706 -3546
rect 85942 -3782 121386 -3546
rect 121622 -3782 121706 -3546
rect 121942 -3782 157386 -3546
rect 157622 -3782 157706 -3546
rect 157942 -3782 193386 -3546
rect 193622 -3782 193706 -3546
rect 193942 -3782 229386 -3546
rect 229622 -3782 229706 -3546
rect 229942 -3782 265386 -3546
rect 265622 -3782 265706 -3546
rect 265942 -3782 301386 -3546
rect 301622 -3782 301706 -3546
rect 301942 -3782 337386 -3546
rect 337622 -3782 337706 -3546
rect 337942 -3782 373386 -3546
rect 373622 -3782 373706 -3546
rect 373942 -3782 409386 -3546
rect 409622 -3782 409706 -3546
rect 409942 -3782 445386 -3546
rect 445622 -3782 445706 -3546
rect 445942 -3782 481386 -3546
rect 481622 -3782 481706 -3546
rect 481942 -3782 517386 -3546
rect 517622 -3782 517706 -3546
rect 517942 -3782 553386 -3546
rect 553622 -3782 553706 -3546
rect 553942 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 17106 -4186
rect 17342 -4422 17426 -4186
rect 17662 -4422 53106 -4186
rect 53342 -4422 53426 -4186
rect 53662 -4422 89106 -4186
rect 89342 -4422 89426 -4186
rect 89662 -4422 125106 -4186
rect 125342 -4422 125426 -4186
rect 125662 -4422 161106 -4186
rect 161342 -4422 161426 -4186
rect 161662 -4422 197106 -4186
rect 197342 -4422 197426 -4186
rect 197662 -4422 233106 -4186
rect 233342 -4422 233426 -4186
rect 233662 -4422 269106 -4186
rect 269342 -4422 269426 -4186
rect 269662 -4422 305106 -4186
rect 305342 -4422 305426 -4186
rect 305662 -4422 341106 -4186
rect 341342 -4422 341426 -4186
rect 341662 -4422 377106 -4186
rect 377342 -4422 377426 -4186
rect 377662 -4422 413106 -4186
rect 413342 -4422 413426 -4186
rect 413662 -4422 449106 -4186
rect 449342 -4422 449426 -4186
rect 449662 -4422 485106 -4186
rect 485342 -4422 485426 -4186
rect 485662 -4422 521106 -4186
rect 521342 -4422 521426 -4186
rect 521662 -4422 557106 -4186
rect 557342 -4422 557426 -4186
rect 557662 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 17106 -4506
rect 17342 -4742 17426 -4506
rect 17662 -4742 53106 -4506
rect 53342 -4742 53426 -4506
rect 53662 -4742 89106 -4506
rect 89342 -4742 89426 -4506
rect 89662 -4742 125106 -4506
rect 125342 -4742 125426 -4506
rect 125662 -4742 161106 -4506
rect 161342 -4742 161426 -4506
rect 161662 -4742 197106 -4506
rect 197342 -4742 197426 -4506
rect 197662 -4742 233106 -4506
rect 233342 -4742 233426 -4506
rect 233662 -4742 269106 -4506
rect 269342 -4742 269426 -4506
rect 269662 -4742 305106 -4506
rect 305342 -4742 305426 -4506
rect 305662 -4742 341106 -4506
rect 341342 -4742 341426 -4506
rect 341662 -4742 377106 -4506
rect 377342 -4742 377426 -4506
rect 377662 -4742 413106 -4506
rect 413342 -4742 413426 -4506
rect 413662 -4742 449106 -4506
rect 449342 -4742 449426 -4506
rect 449662 -4742 485106 -4506
rect 485342 -4742 485426 -4506
rect 485662 -4742 521106 -4506
rect 521342 -4742 521426 -4506
rect 521662 -4742 557106 -4506
rect 557342 -4742 557426 -4506
rect 557662 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20826 -5146
rect 21062 -5382 21146 -5146
rect 21382 -5382 56826 -5146
rect 57062 -5382 57146 -5146
rect 57382 -5382 92826 -5146
rect 93062 -5382 93146 -5146
rect 93382 -5382 128826 -5146
rect 129062 -5382 129146 -5146
rect 129382 -5382 164826 -5146
rect 165062 -5382 165146 -5146
rect 165382 -5382 200826 -5146
rect 201062 -5382 201146 -5146
rect 201382 -5382 236826 -5146
rect 237062 -5382 237146 -5146
rect 237382 -5382 272826 -5146
rect 273062 -5382 273146 -5146
rect 273382 -5382 308826 -5146
rect 309062 -5382 309146 -5146
rect 309382 -5382 344826 -5146
rect 345062 -5382 345146 -5146
rect 345382 -5382 380826 -5146
rect 381062 -5382 381146 -5146
rect 381382 -5382 416826 -5146
rect 417062 -5382 417146 -5146
rect 417382 -5382 452826 -5146
rect 453062 -5382 453146 -5146
rect 453382 -5382 488826 -5146
rect 489062 -5382 489146 -5146
rect 489382 -5382 524826 -5146
rect 525062 -5382 525146 -5146
rect 525382 -5382 560826 -5146
rect 561062 -5382 561146 -5146
rect 561382 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20826 -5466
rect 21062 -5702 21146 -5466
rect 21382 -5702 56826 -5466
rect 57062 -5702 57146 -5466
rect 57382 -5702 92826 -5466
rect 93062 -5702 93146 -5466
rect 93382 -5702 128826 -5466
rect 129062 -5702 129146 -5466
rect 129382 -5702 164826 -5466
rect 165062 -5702 165146 -5466
rect 165382 -5702 200826 -5466
rect 201062 -5702 201146 -5466
rect 201382 -5702 236826 -5466
rect 237062 -5702 237146 -5466
rect 237382 -5702 272826 -5466
rect 273062 -5702 273146 -5466
rect 273382 -5702 308826 -5466
rect 309062 -5702 309146 -5466
rect 309382 -5702 344826 -5466
rect 345062 -5702 345146 -5466
rect 345382 -5702 380826 -5466
rect 381062 -5702 381146 -5466
rect 381382 -5702 416826 -5466
rect 417062 -5702 417146 -5466
rect 417382 -5702 452826 -5466
rect 453062 -5702 453146 -5466
rect 453382 -5702 488826 -5466
rect 489062 -5702 489146 -5466
rect 489382 -5702 524826 -5466
rect 525062 -5702 525146 -5466
rect 525382 -5702 560826 -5466
rect 561062 -5702 561146 -5466
rect 561382 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24546 -6106
rect 24782 -6342 24866 -6106
rect 25102 -6342 60546 -6106
rect 60782 -6342 60866 -6106
rect 61102 -6342 96546 -6106
rect 96782 -6342 96866 -6106
rect 97102 -6342 132546 -6106
rect 132782 -6342 132866 -6106
rect 133102 -6342 168546 -6106
rect 168782 -6342 168866 -6106
rect 169102 -6342 204546 -6106
rect 204782 -6342 204866 -6106
rect 205102 -6342 240546 -6106
rect 240782 -6342 240866 -6106
rect 241102 -6342 276546 -6106
rect 276782 -6342 276866 -6106
rect 277102 -6342 312546 -6106
rect 312782 -6342 312866 -6106
rect 313102 -6342 348546 -6106
rect 348782 -6342 348866 -6106
rect 349102 -6342 384546 -6106
rect 384782 -6342 384866 -6106
rect 385102 -6342 420546 -6106
rect 420782 -6342 420866 -6106
rect 421102 -6342 456546 -6106
rect 456782 -6342 456866 -6106
rect 457102 -6342 492546 -6106
rect 492782 -6342 492866 -6106
rect 493102 -6342 528546 -6106
rect 528782 -6342 528866 -6106
rect 529102 -6342 564546 -6106
rect 564782 -6342 564866 -6106
rect 565102 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24546 -6426
rect 24782 -6662 24866 -6426
rect 25102 -6662 60546 -6426
rect 60782 -6662 60866 -6426
rect 61102 -6662 96546 -6426
rect 96782 -6662 96866 -6426
rect 97102 -6662 132546 -6426
rect 132782 -6662 132866 -6426
rect 133102 -6662 168546 -6426
rect 168782 -6662 168866 -6426
rect 169102 -6662 204546 -6426
rect 204782 -6662 204866 -6426
rect 205102 -6662 240546 -6426
rect 240782 -6662 240866 -6426
rect 241102 -6662 276546 -6426
rect 276782 -6662 276866 -6426
rect 277102 -6662 312546 -6426
rect 312782 -6662 312866 -6426
rect 313102 -6662 348546 -6426
rect 348782 -6662 348866 -6426
rect 349102 -6662 384546 -6426
rect 384782 -6662 384866 -6426
rect 385102 -6662 420546 -6426
rect 420782 -6662 420866 -6426
rect 421102 -6662 456546 -6426
rect 456782 -6662 456866 -6426
rect 457102 -6662 492546 -6426
rect 492782 -6662 492866 -6426
rect 493102 -6662 528546 -6426
rect 528782 -6662 528866 -6426
rect 529102 -6662 564546 -6426
rect 564782 -6662 564866 -6426
rect 565102 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 28266 -7066
rect 28502 -7302 28586 -7066
rect 28822 -7302 64266 -7066
rect 64502 -7302 64586 -7066
rect 64822 -7302 100266 -7066
rect 100502 -7302 100586 -7066
rect 100822 -7302 136266 -7066
rect 136502 -7302 136586 -7066
rect 136822 -7302 172266 -7066
rect 172502 -7302 172586 -7066
rect 172822 -7302 208266 -7066
rect 208502 -7302 208586 -7066
rect 208822 -7302 244266 -7066
rect 244502 -7302 244586 -7066
rect 244822 -7302 280266 -7066
rect 280502 -7302 280586 -7066
rect 280822 -7302 316266 -7066
rect 316502 -7302 316586 -7066
rect 316822 -7302 352266 -7066
rect 352502 -7302 352586 -7066
rect 352822 -7302 388266 -7066
rect 388502 -7302 388586 -7066
rect 388822 -7302 424266 -7066
rect 424502 -7302 424586 -7066
rect 424822 -7302 460266 -7066
rect 460502 -7302 460586 -7066
rect 460822 -7302 496266 -7066
rect 496502 -7302 496586 -7066
rect 496822 -7302 532266 -7066
rect 532502 -7302 532586 -7066
rect 532822 -7302 568266 -7066
rect 568502 -7302 568586 -7066
rect 568822 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 28266 -7386
rect 28502 -7622 28586 -7386
rect 28822 -7622 64266 -7386
rect 64502 -7622 64586 -7386
rect 64822 -7622 100266 -7386
rect 100502 -7622 100586 -7386
rect 100822 -7622 136266 -7386
rect 136502 -7622 136586 -7386
rect 136822 -7622 172266 -7386
rect 172502 -7622 172586 -7386
rect 172822 -7622 208266 -7386
rect 208502 -7622 208586 -7386
rect 208822 -7622 244266 -7386
rect 244502 -7622 244586 -7386
rect 244822 -7622 280266 -7386
rect 280502 -7622 280586 -7386
rect 280822 -7622 316266 -7386
rect 316502 -7622 316586 -7386
rect 316822 -7622 352266 -7386
rect 352502 -7622 352586 -7386
rect 352822 -7622 388266 -7386
rect 388502 -7622 388586 -7386
rect 388822 -7622 424266 -7386
rect 424502 -7622 424586 -7386
rect 424822 -7622 460266 -7386
rect 460502 -7622 460586 -7386
rect 460822 -7622 496266 -7386
rect 496502 -7622 496586 -7386
rect 496822 -7622 532266 -7386
rect 532502 -7622 532586 -7386
rect 532822 -7622 568266 -7386
rect 568502 -7622 568586 -7386
rect 568822 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use egd_top_wrapper  egd_top_wrapper
timestamp 0
transform 1 0 400000 0 1 80000
box 0 0 52610 53360
use R4_butter  R4_butter
timestamp 0
transform 1 0 300000 0 1 80000
box 1066 0 36400 38800
use wb_buttons_leds  wb_buttons_leds
timestamp 0
transform 1 0 80000 0 1 80000
box 1066 0 110000 110000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 2194 -7654 2814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 38194 -7654 38814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 74194 -7654 74814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 110194 -7654 110814 81159 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 110194 188457 110814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 146194 -7654 146814 81159 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 146194 188457 146814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 182194 -7654 182814 81159 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 182194 188457 182814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 218194 -7654 218814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 254194 -7654 254814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 290194 -7654 290814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 326194 -7654 326814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 362194 -7654 362814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 398194 -7654 398814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 434194 -7654 434814 79988 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 434194 135500 434814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 470194 -7654 470814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 506194 -7654 506814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 542194 -7654 542814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 578194 -7654 578814 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 3266 592650 3886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 39266 592650 39886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 75266 592650 75886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 111266 592650 111886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 147266 592650 147886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 183266 592650 183886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 219266 592650 219886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 255266 592650 255886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 291266 592650 291886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 327266 592650 327886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 363266 592650 363886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 399266 592650 399886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 435266 592650 435886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 471266 592650 471886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 507266 592650 507886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 543266 592650 543886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 579266 592650 579886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 615266 592650 615886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 651266 592650 651886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 687266 592650 687886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9634 -7654 10254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45634 -7654 46254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81634 -7654 82254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117634 -7654 118254 81159 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117634 188457 118254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153634 -7654 154254 81159 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153634 188457 154254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189634 -7654 190254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225634 -7654 226254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261634 -7654 262254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297634 -7654 298254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333634 -7654 334254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369634 -7654 370254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405634 -7654 406254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441634 -7654 442254 81159 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441634 133649 442254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477634 -7654 478254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513634 -7654 514254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549634 -7654 550254 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10706 592650 11326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46706 592650 47326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82706 592650 83326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118706 592650 119326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154706 592650 155326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190706 592650 191326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226706 592650 227326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262706 592650 263326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298706 592650 299326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334706 592650 335326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370706 592650 371326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406706 592650 407326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442706 592650 443326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478706 592650 479326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514706 592650 515326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550706 592650 551326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586706 592650 587326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622706 592650 623326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658706 592650 659326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694706 592650 695326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 17074 -7654 17694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 53074 -7654 53694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 89074 -7654 89694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 125074 -7654 125694 81159 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 125074 188457 125694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 161074 -7654 161694 79988 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 161074 189900 161694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 197074 -7654 197694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 233074 -7654 233694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 269074 -7654 269694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 305074 -7654 305694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 341074 -7654 341694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 377074 -7654 377694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 413074 -7654 413694 81159 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 413074 133649 413694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 449074 -7654 449694 81159 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 449074 133649 449694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 485074 -7654 485694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 521074 -7654 521694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 557074 -7654 557694 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 18146 592650 18766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 54146 592650 54766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 90146 592650 90766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 126146 592650 126766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 162146 592650 162766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 198146 592650 198766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 234146 592650 234766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 270146 592650 270766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 306146 592650 306766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 342146 592650 342766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 378146 592650 378766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 414146 592650 414766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 450146 592650 450766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 486146 592650 486766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 522146 592650 522766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 558146 592650 558766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 594146 592650 594766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 630146 592650 630766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 666146 592650 666766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24514 -7654 25134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60514 -7654 61134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96514 -7654 97134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132514 -7654 133134 81159 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132514 188457 133134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168514 -7654 169134 81159 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168514 188457 169134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204514 -7654 205134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240514 -7654 241134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276514 -7654 277134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312514 -7654 313134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348514 -7654 349134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384514 -7654 385134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420514 -7654 421134 81159 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420514 133586 421134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456514 -7654 457134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492514 -7654 493134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528514 -7654 529134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564514 -7654 565134 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25586 592650 26206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61586 592650 62206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97586 592650 98206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133586 592650 134206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169586 592650 170206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205586 592650 206206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241586 592650 242206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277586 592650 278206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313586 592650 314206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349586 592650 350206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385586 592650 386206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421586 592650 422206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457586 592650 458206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493586 592650 494206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529586 592650 530206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565586 592650 566206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601586 592650 602206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637586 592650 638206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673586 592650 674206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20794 -7654 21414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56794 -7654 57414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92794 -7654 93414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128794 -7654 129414 81159 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128794 188457 129414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164794 -7654 165414 81159 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164794 188457 165414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200794 -7654 201414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236794 -7654 237414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272794 -7654 273414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308794 -7654 309414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344794 -7654 345414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380794 -7654 381414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416794 -7654 417414 81159 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416794 133649 417414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452794 -7654 453414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488794 -7654 489414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524794 -7654 525414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560794 -7654 561414 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21866 592650 22486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57866 592650 58486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93866 592650 94486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129866 592650 130486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165866 592650 166486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201866 592650 202486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237866 592650 238486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273866 592650 274486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309866 592650 310486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345866 592650 346486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381866 592650 382486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417866 592650 418486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453866 592650 454486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489866 592650 490486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525866 592650 526486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561866 592650 562486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597866 592650 598486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633866 592650 634486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669866 592650 670486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 28234 -7654 28854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 64234 -7654 64854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 100234 -7654 100854 81159 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 100234 188457 100854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 136234 -7654 136854 81159 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 136234 188457 136854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 172234 -7654 172854 81159 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 172234 188457 172854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 208234 -7654 208854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 244234 -7654 244854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 280234 -7654 280854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 316234 -7654 316854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 352234 -7654 352854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 388234 -7654 388854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 424234 -7654 424854 81159 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 424234 133649 424854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 460234 -7654 460854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 496234 -7654 496854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 532234 -7654 532854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 568234 -7654 568854 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 29306 592650 29926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 65306 592650 65926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 101306 592650 101926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 137306 592650 137926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 173306 592650 173926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 209306 592650 209926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 245306 592650 245926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 281306 592650 281926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 317306 592650 317926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 353306 592650 353926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 389306 592650 389926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 425306 592650 425926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 461306 592650 461926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 497306 592650 497926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 533306 592650 533926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 569306 592650 569926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 605306 592650 605926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 641306 592650 641926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 677306 592650 677926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5914 -7654 6534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41914 -7654 42534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77914 -7654 78534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113914 -7654 114534 81159 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113914 188457 114534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149914 -7654 150534 81159 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149914 188457 150534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185914 -7654 186534 81159 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185914 188457 186534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221914 -7654 222534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257914 -7654 258534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293914 -7654 294534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329914 -7654 330534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365914 -7654 366534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401914 -7654 402534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437914 -7654 438534 81159 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437914 133649 438534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473914 -7654 474534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509914 -7654 510534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545914 -7654 546534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581914 -7654 582534 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6986 592650 7606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42986 592650 43606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78986 592650 79606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114986 592650 115606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150986 592650 151606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186986 592650 187606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222986 592650 223606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258986 592650 259606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294986 592650 295606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330986 592650 331606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366986 592650 367606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402986 592650 403606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438986 592650 439606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474986 592650 475606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510986 592650 511606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546986 592650 547606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582986 592650 583606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618986 592650 619606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654986 592650 655606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690986 592650 691606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 13354 -7654 13974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 49354 -7654 49974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 85354 -7654 85974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 121354 -7654 121974 81159 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 121354 188457 121974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 157354 -7654 157974 81159 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 157354 188457 157974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 193354 -7654 193974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 229354 -7654 229974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 265354 -7654 265974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 301354 -7654 301974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 337354 -7654 337974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 373354 -7654 373974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 409354 -7654 409974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 445354 -7654 445974 81159 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 445354 133649 445974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 481354 -7654 481974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 517354 -7654 517974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 553354 -7654 553974 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14426 592650 15046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50426 592650 51046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86426 592650 87046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122426 592650 123046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158426 592650 159046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194426 592650 195046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230426 592650 231046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266426 592650 267046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302426 592650 303046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338426 592650 339046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374426 592650 375046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410426 592650 411046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446426 592650 447046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482426 592650 483046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518426 592650 519046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554426 592650 555046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590426 592650 591046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626426 592650 627046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662426 592650 663046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698426 592650 699046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
