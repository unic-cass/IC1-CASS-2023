magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 10 76 554 730
<< nmoslvt >>
rect 204 102 254 704
rect 310 102 360 704
<< ndiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 254 692 310 704
rect 254 658 265 692
rect 299 658 310 692
rect 254 624 310 658
rect 254 590 265 624
rect 299 590 310 624
rect 254 556 310 590
rect 254 522 265 556
rect 299 522 310 556
rect 254 488 310 522
rect 254 454 265 488
rect 299 454 310 488
rect 254 420 310 454
rect 254 386 265 420
rect 299 386 310 420
rect 254 352 310 386
rect 254 318 265 352
rect 299 318 310 352
rect 254 284 310 318
rect 254 250 265 284
rect 299 250 310 284
rect 254 216 310 250
rect 254 182 265 216
rect 299 182 310 216
rect 254 148 310 182
rect 254 114 265 148
rect 299 114 310 148
rect 254 102 310 114
rect 360 692 416 704
rect 360 658 371 692
rect 405 658 416 692
rect 360 624 416 658
rect 360 590 371 624
rect 405 590 416 624
rect 360 556 416 590
rect 360 522 371 556
rect 405 522 416 556
rect 360 488 416 522
rect 360 454 371 488
rect 405 454 416 488
rect 360 420 416 454
rect 360 386 371 420
rect 405 386 416 420
rect 360 352 416 386
rect 360 318 371 352
rect 405 318 416 352
rect 360 284 416 318
rect 360 250 371 284
rect 405 250 416 284
rect 360 216 416 250
rect 360 182 371 216
rect 405 182 416 216
rect 360 148 416 182
rect 360 114 371 148
rect 405 114 416 148
rect 360 102 416 114
<< ndiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 265 658 299 692
rect 265 590 299 624
rect 265 522 299 556
rect 265 454 299 488
rect 265 386 299 420
rect 265 318 299 352
rect 265 250 299 284
rect 265 182 299 216
rect 265 114 299 148
rect 371 658 405 692
rect 371 590 405 624
rect 371 522 405 556
rect 371 454 405 488
rect 371 386 405 420
rect 371 318 405 352
rect 371 250 405 284
rect 371 182 405 216
rect 371 114 405 148
<< psubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 470 658 528 704
rect 470 624 482 658
rect 516 624 528 658
rect 470 590 528 624
rect 470 556 482 590
rect 516 556 528 590
rect 470 522 528 556
rect 470 488 482 522
rect 516 488 528 522
rect 470 454 528 488
rect 470 420 482 454
rect 516 420 528 454
rect 470 386 528 420
rect 470 352 482 386
rect 516 352 528 386
rect 470 318 528 352
rect 470 284 482 318
rect 516 284 528 318
rect 470 250 528 284
rect 470 216 482 250
rect 516 216 528 250
rect 470 182 528 216
rect 470 148 482 182
rect 516 148 528 182
rect 470 102 528 148
<< psubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 482 624 516 658
rect 482 556 516 590
rect 482 488 516 522
rect 482 420 516 454
rect 482 352 516 386
rect 482 284 516 318
rect 482 216 516 250
rect 482 148 516 182
<< poly >>
rect 181 776 383 796
rect 181 742 197 776
rect 231 742 265 776
rect 299 742 333 776
rect 367 742 383 776
rect 181 726 383 742
rect 204 704 254 726
rect 310 704 360 726
rect 204 80 254 102
rect 310 80 360 102
rect 181 64 383 80
rect 181 30 197 64
rect 231 30 265 64
rect 299 30 333 64
rect 367 30 383 64
rect 181 10 383 30
<< polycont >>
rect 197 742 231 776
rect 265 742 299 776
rect 333 742 367 776
rect 197 30 231 64
rect 265 30 299 64
rect 333 30 367 64
<< locali >>
rect 181 742 193 776
rect 231 742 265 776
rect 299 742 333 776
rect 371 742 383 776
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 265 692 299 708
rect 265 624 299 638
rect 265 556 299 566
rect 265 488 299 494
rect 265 420 299 422
rect 265 384 299 386
rect 265 312 299 318
rect 265 240 299 250
rect 265 168 299 182
rect 265 98 299 114
rect 371 692 405 708
rect 371 624 405 638
rect 371 556 405 566
rect 371 488 405 494
rect 371 420 405 422
rect 371 384 405 386
rect 371 312 405 318
rect 371 240 405 250
rect 371 168 405 182
rect 482 672 516 674
rect 482 600 516 624
rect 482 528 516 556
rect 482 456 516 488
rect 482 386 516 420
rect 482 318 516 350
rect 482 250 516 278
rect 482 182 516 206
rect 482 132 516 134
rect 371 98 405 114
rect 181 30 193 64
rect 231 30 265 64
rect 299 30 333 64
rect 371 30 383 64
<< viali >>
rect 193 742 197 776
rect 197 742 227 776
rect 265 742 299 776
rect 337 742 367 776
rect 367 742 371 776
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 265 658 299 672
rect 265 638 299 658
rect 265 590 299 600
rect 265 566 299 590
rect 265 522 299 528
rect 265 494 299 522
rect 265 454 299 456
rect 265 422 299 454
rect 265 352 299 384
rect 265 350 299 352
rect 265 284 299 312
rect 265 278 299 284
rect 265 216 299 240
rect 265 206 299 216
rect 265 148 299 168
rect 265 134 299 148
rect 371 658 405 672
rect 371 638 405 658
rect 371 590 405 600
rect 371 566 405 590
rect 371 522 405 528
rect 371 494 405 522
rect 371 454 405 456
rect 371 422 405 454
rect 371 352 405 384
rect 371 350 405 352
rect 371 284 405 312
rect 371 278 405 284
rect 371 216 405 240
rect 371 206 405 216
rect 371 148 405 168
rect 371 134 405 148
rect 482 658 516 672
rect 482 638 516 658
rect 482 590 516 600
rect 482 566 516 590
rect 482 522 516 528
rect 482 494 516 522
rect 482 454 516 456
rect 482 422 516 454
rect 482 352 516 384
rect 482 350 516 352
rect 482 284 516 312
rect 482 278 516 284
rect 482 216 516 240
rect 482 206 516 216
rect 482 148 516 168
rect 482 134 516 148
rect 193 30 197 64
rect 197 30 227 64
rect 265 30 299 64
rect 337 30 367 64
rect 367 30 371 64
<< metal1 >>
rect 181 776 383 796
rect 181 742 193 776
rect 227 742 265 776
rect 299 742 337 776
rect 371 742 383 776
rect 181 730 383 742
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 256 678 308 684
rect 256 614 308 626
rect 256 550 308 562
rect 256 494 265 498
rect 299 494 308 498
rect 256 486 308 494
rect 256 422 265 434
rect 299 422 308 434
rect 256 384 308 422
rect 256 350 265 384
rect 299 350 308 384
rect 256 312 308 350
rect 256 278 265 312
rect 299 278 308 312
rect 256 240 308 278
rect 256 206 265 240
rect 299 206 308 240
rect 256 168 308 206
rect 256 134 265 168
rect 299 134 308 168
rect 256 122 308 134
rect 362 672 414 684
rect 362 638 371 672
rect 405 638 414 672
rect 362 600 414 638
rect 362 566 371 600
rect 405 566 414 600
rect 362 528 414 566
rect 362 494 371 528
rect 405 494 414 528
rect 362 456 414 494
rect 362 422 371 456
rect 405 422 414 456
rect 362 384 414 422
rect 362 372 371 384
rect 405 372 414 384
rect 362 312 414 320
rect 362 308 371 312
rect 405 308 414 312
rect 362 244 414 256
rect 362 180 414 192
rect 362 122 414 128
rect 470 672 528 684
rect 470 638 482 672
rect 516 638 528 672
rect 470 600 528 638
rect 470 566 482 600
rect 516 566 528 600
rect 470 528 528 566
rect 470 494 482 528
rect 516 494 528 528
rect 470 456 528 494
rect 470 422 482 456
rect 516 422 528 456
rect 470 384 528 422
rect 470 350 482 384
rect 516 350 528 384
rect 470 312 528 350
rect 470 278 482 312
rect 516 278 528 312
rect 470 240 528 278
rect 470 206 482 240
rect 516 206 528 240
rect 470 168 528 206
rect 470 134 482 168
rect 516 134 528 168
rect 470 122 528 134
rect 181 64 383 76
rect 181 30 193 64
rect 227 30 265 64
rect 299 30 337 64
rect 371 30 383 64
rect 181 10 383 30
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 256 672 308 678
rect 256 638 265 672
rect 265 638 299 672
rect 299 638 308 672
rect 256 626 308 638
rect 256 600 308 614
rect 256 566 265 600
rect 265 566 299 600
rect 299 566 308 600
rect 256 562 308 566
rect 256 528 308 550
rect 256 498 265 528
rect 265 498 299 528
rect 299 498 308 528
rect 256 456 308 486
rect 256 434 265 456
rect 265 434 299 456
rect 299 434 308 456
rect 362 350 371 372
rect 371 350 405 372
rect 405 350 414 372
rect 362 320 414 350
rect 362 278 371 308
rect 371 278 405 308
rect 405 278 414 308
rect 362 256 414 278
rect 362 240 414 244
rect 362 206 371 240
rect 371 206 405 240
rect 405 206 414 240
rect 362 192 414 206
rect 362 168 414 180
rect 362 134 371 168
rect 371 134 405 168
rect 405 134 414 168
rect 362 128 414 134
<< metal2 >>
rect 10 678 554 684
rect 10 626 256 678
rect 308 626 554 678
rect 10 614 554 626
rect 10 562 256 614
rect 308 562 554 614
rect 10 550 554 562
rect 10 498 256 550
rect 308 498 554 550
rect 10 486 554 498
rect 10 434 256 486
rect 308 434 554 486
rect 10 428 554 434
rect 10 372 554 378
rect 10 320 150 372
rect 202 320 362 372
rect 414 320 554 372
rect 10 308 554 320
rect 10 256 150 308
rect 202 256 362 308
rect 414 256 554 308
rect 10 244 554 256
rect 10 192 150 244
rect 202 192 362 244
rect 414 192 554 244
rect 10 180 554 192
rect 10 128 150 180
rect 202 128 362 180
rect 414 128 554 180
rect 10 122 554 128
<< labels >>
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
port 2 nsew
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
port 3 nsew
flabel metal1 s 181 730 383 796 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 181 10 383 76 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 470 122 528 138 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
<< properties >>
string GDS_END 3453912
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3442984
<< end >>
