magic
tech sky130A
magscale 1 2
timestamp 1698801821
<< nwell >>
rect 1066 36165 35274 36486
rect 1066 35077 35274 35643
rect 1066 33989 35274 34555
rect 1066 32901 35274 33467
rect 1066 31813 35274 32379
rect 1066 30725 35274 31291
rect 1066 29637 35274 30203
rect 1066 28549 35274 29115
rect 1066 27461 35274 28027
rect 1066 26373 35274 26939
rect 1066 25285 35274 25851
rect 1066 24197 35274 24763
rect 1066 23109 35274 23675
rect 1066 22021 35274 22587
rect 1066 20933 35274 21499
rect 1066 19845 35274 20411
rect 1066 18757 35274 19323
rect 1066 17669 35274 18235
rect 1066 16581 35274 17147
rect 1066 15493 35274 16059
rect 1066 14405 35274 14971
rect 1066 13317 35274 13883
rect 1066 12229 35274 12795
rect 1066 11141 35274 11707
rect 1066 10053 35274 10619
rect 1066 8965 35274 9531
rect 1066 7877 35274 8443
rect 1066 6789 35274 7355
rect 1066 5701 35274 6267
rect 1066 4613 35274 5179
rect 1066 3525 35274 4091
rect 1066 2437 35274 3003
<< obsli1 >>
rect 1104 2159 35236 36465
<< obsm1 >>
rect 1104 2128 35866 36496
<< metal2 >>
rect 4526 38000 4582 38800
rect 13634 38000 13690 38800
rect 22742 38000 22798 38800
rect 31850 38000 31906 38800
rect 2410 0 2466 800
rect 6918 0 6974 800
rect 11426 0 11482 800
rect 15934 0 15990 800
rect 20442 0 20498 800
rect 24950 0 25006 800
rect 29458 0 29514 800
rect 33966 0 34022 800
<< obsm2 >>
rect 2412 37944 4470 38162
rect 4638 37944 13578 38162
rect 13746 37944 22686 38162
rect 22854 37944 31794 38162
rect 31962 37944 35860 38162
rect 2412 856 35860 37944
rect 2522 800 6862 856
rect 7030 800 11370 856
rect 11538 800 15878 856
rect 16046 800 20386 856
rect 20554 800 24894 856
rect 25062 800 29402 856
rect 29570 800 33910 856
rect 34078 800 35860 856
<< metal3 >>
rect 35600 37408 36400 37528
rect 35600 36456 36400 36576
rect 35600 35504 36400 35624
rect 35600 34552 36400 34672
rect 35600 33600 36400 33720
rect 35600 32648 36400 32768
rect 35600 31696 36400 31816
rect 35600 30744 36400 30864
rect 35600 29792 36400 29912
rect 35600 28840 36400 28960
rect 35600 27888 36400 28008
rect 35600 26936 36400 27056
rect 35600 25984 36400 26104
rect 35600 25032 36400 25152
rect 35600 24080 36400 24200
rect 35600 23128 36400 23248
rect 35600 22176 36400 22296
rect 35600 21224 36400 21344
rect 35600 20272 36400 20392
rect 35600 19320 36400 19440
rect 35600 18368 36400 18488
rect 35600 17416 36400 17536
rect 35600 16464 36400 16584
rect 35600 15512 36400 15632
rect 35600 14560 36400 14680
rect 35600 13608 36400 13728
rect 35600 12656 36400 12776
rect 35600 11704 36400 11824
rect 35600 10752 36400 10872
rect 35600 9800 36400 9920
rect 35600 8848 36400 8968
rect 35600 7896 36400 8016
rect 35600 6944 36400 7064
rect 35600 5992 36400 6112
rect 35600 5040 36400 5160
rect 35600 4088 36400 4208
rect 35600 3136 36400 3256
rect 35600 2184 36400 2304
rect 35600 1232 36400 1352
<< obsm3 >>
rect 4210 37328 35520 37501
rect 4210 36656 35600 37328
rect 4210 36376 35520 36656
rect 4210 35704 35600 36376
rect 4210 35424 35520 35704
rect 4210 34752 35600 35424
rect 4210 34472 35520 34752
rect 4210 33800 35600 34472
rect 4210 33520 35520 33800
rect 4210 32848 35600 33520
rect 4210 32568 35520 32848
rect 4210 31896 35600 32568
rect 4210 31616 35520 31896
rect 4210 30944 35600 31616
rect 4210 30664 35520 30944
rect 4210 29992 35600 30664
rect 4210 29712 35520 29992
rect 4210 29040 35600 29712
rect 4210 28760 35520 29040
rect 4210 28088 35600 28760
rect 4210 27808 35520 28088
rect 4210 27136 35600 27808
rect 4210 26856 35520 27136
rect 4210 26184 35600 26856
rect 4210 25904 35520 26184
rect 4210 25232 35600 25904
rect 4210 24952 35520 25232
rect 4210 24280 35600 24952
rect 4210 24000 35520 24280
rect 4210 23328 35600 24000
rect 4210 23048 35520 23328
rect 4210 22376 35600 23048
rect 4210 22096 35520 22376
rect 4210 21424 35600 22096
rect 4210 21144 35520 21424
rect 4210 20472 35600 21144
rect 4210 20192 35520 20472
rect 4210 19520 35600 20192
rect 4210 19240 35520 19520
rect 4210 18568 35600 19240
rect 4210 18288 35520 18568
rect 4210 17616 35600 18288
rect 4210 17336 35520 17616
rect 4210 16664 35600 17336
rect 4210 16384 35520 16664
rect 4210 15712 35600 16384
rect 4210 15432 35520 15712
rect 4210 14760 35600 15432
rect 4210 14480 35520 14760
rect 4210 13808 35600 14480
rect 4210 13528 35520 13808
rect 4210 12856 35600 13528
rect 4210 12576 35520 12856
rect 4210 11904 35600 12576
rect 4210 11624 35520 11904
rect 4210 10952 35600 11624
rect 4210 10672 35520 10952
rect 4210 10000 35600 10672
rect 4210 9720 35520 10000
rect 4210 9048 35600 9720
rect 4210 8768 35520 9048
rect 4210 8096 35600 8768
rect 4210 7816 35520 8096
rect 4210 7144 35600 7816
rect 4210 6864 35520 7144
rect 4210 6192 35600 6864
rect 4210 5912 35520 6192
rect 4210 5240 35600 5912
rect 4210 4960 35520 5240
rect 4210 4288 35600 4960
rect 4210 4008 35520 4288
rect 4210 3336 35600 4008
rect 4210 3056 35520 3336
rect 4210 2384 35600 3056
rect 4210 2104 35520 2384
rect 4210 1432 35600 2104
rect 4210 1259 35520 1432
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< labels >>
rlabel metal3 s 35600 9800 36400 9920 6 Xio[0]
port 1 nsew signal output
rlabel metal3 s 35600 19320 36400 19440 6 Xio[1]
port 2 nsew signal output
rlabel metal3 s 35600 28840 36400 28960 6 Xio[2]
port 3 nsew signal output
rlabel metal3 s 35600 37408 36400 37528 6 Xio[3]
port 4 nsew signal output
rlabel metal3 s 35600 8848 36400 8968 6 Xro[0]
port 5 nsew signal output
rlabel metal3 s 35600 18368 36400 18488 6 Xro[1]
port 6 nsew signal output
rlabel metal3 s 35600 27888 36400 28008 6 Xro[2]
port 7 nsew signal output
rlabel metal3 s 35600 36456 36400 36576 6 Xro[3]
port 8 nsew signal output
rlabel metal2 s 4526 38000 4582 38800 6 c1
port 9 nsew signal input
rlabel metal2 s 13634 38000 13690 38800 6 c2
port 10 nsew signal input
rlabel metal2 s 22742 38000 22798 38800 6 c3
port 11 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 la_oenb[0]
port 12 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 la_oenb[1]
port 13 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 la_oenb[2]
port 14 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 la_oenb[3]
port 15 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 la_oenb[4]
port 16 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_oenb[5]
port 17 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_oenb[6]
port 18 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_oenb[7]
port 19 nsew signal output
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 20 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 20 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 21 nsew ground bidirectional
rlabel metal3 s 35600 2184 36400 2304 6 xi0[0]
port 22 nsew signal input
rlabel metal3 s 35600 11704 36400 11824 6 xi0[1]
port 23 nsew signal input
rlabel metal3 s 35600 21224 36400 21344 6 xi0[2]
port 24 nsew signal input
rlabel metal3 s 35600 30744 36400 30864 6 xi0[3]
port 25 nsew signal input
rlabel metal3 s 35600 4088 36400 4208 6 xi1[0]
port 26 nsew signal input
rlabel metal3 s 35600 13608 36400 13728 6 xi1[1]
port 27 nsew signal input
rlabel metal3 s 35600 23128 36400 23248 6 xi1[2]
port 28 nsew signal input
rlabel metal3 s 35600 32648 36400 32768 6 xi1[3]
port 29 nsew signal input
rlabel metal3 s 35600 5992 36400 6112 6 xi2[0]
port 30 nsew signal input
rlabel metal3 s 35600 15512 36400 15632 6 xi2[1]
port 31 nsew signal input
rlabel metal3 s 35600 25032 36400 25152 6 xi2[2]
port 32 nsew signal input
rlabel metal3 s 35600 34552 36400 34672 6 xi2[3]
port 33 nsew signal input
rlabel metal3 s 35600 7896 36400 8016 6 xi3[0]
port 34 nsew signal input
rlabel metal3 s 35600 17416 36400 17536 6 xi3[1]
port 35 nsew signal input
rlabel metal3 s 35600 26936 36400 27056 6 xi3[2]
port 36 nsew signal input
rlabel metal2 s 31850 38000 31906 38800 6 xi3[3]
port 37 nsew signal input
rlabel metal3 s 35600 1232 36400 1352 6 xr0[0]
port 38 nsew signal input
rlabel metal3 s 35600 10752 36400 10872 6 xr0[1]
port 39 nsew signal input
rlabel metal3 s 35600 20272 36400 20392 6 xr0[2]
port 40 nsew signal input
rlabel metal3 s 35600 29792 36400 29912 6 xr0[3]
port 41 nsew signal input
rlabel metal3 s 35600 3136 36400 3256 6 xr1[0]
port 42 nsew signal input
rlabel metal3 s 35600 12656 36400 12776 6 xr1[1]
port 43 nsew signal input
rlabel metal3 s 35600 22176 36400 22296 6 xr1[2]
port 44 nsew signal input
rlabel metal3 s 35600 31696 36400 31816 6 xr1[3]
port 45 nsew signal input
rlabel metal3 s 35600 5040 36400 5160 6 xr2[0]
port 46 nsew signal input
rlabel metal3 s 35600 14560 36400 14680 6 xr2[1]
port 47 nsew signal input
rlabel metal3 s 35600 24080 36400 24200 6 xr2[2]
port 48 nsew signal input
rlabel metal3 s 35600 33600 36400 33720 6 xr2[3]
port 49 nsew signal input
rlabel metal3 s 35600 6944 36400 7064 6 xr3[0]
port 50 nsew signal input
rlabel metal3 s 35600 16464 36400 16584 6 xr3[1]
port 51 nsew signal input
rlabel metal3 s 35600 25984 36400 26104 6 xr3[2]
port 52 nsew signal input
rlabel metal3 s 35600 35504 36400 35624 6 xr3[3]
port 53 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36400 38800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 435208
string GDS_FILE /home/rodrigowue/IC1-V2/openlane/R4_butter/runs/23_10_31_22_22/results/signoff/R4_butter.magic.gds
string GDS_START 44362
<< end >>

