magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 3074 582
<< pwell >>
rect 2398 201 3035 203
rect 1241 157 1695 201
rect 2016 157 3035 201
rect 1 21 3035 157
rect 29 -17 63 21
<< locali >>
rect 17 195 87 325
rect 283 205 339 337
rect 387 219 431 339
rect 387 153 467 219
rect 765 265 805 475
rect 387 69 429 153
rect 2516 326 2566 493
rect 2318 219 2414 265
rect 2532 143 2566 326
rect 2883 289 2933 493
rect 2516 51 2566 143
rect 2892 165 2933 289
rect 2883 51 2933 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 34 393 69 493
rect 103 427 169 527
rect 34 359 167 393
rect 121 161 167 359
rect 34 127 167 161
rect 34 69 69 127
rect 103 17 169 93
rect 203 69 247 493
rect 286 377 357 527
rect 443 375 515 477
rect 579 381 613 493
rect 659 443 728 527
rect 481 281 515 375
rect 549 349 613 381
rect 549 315 729 349
rect 481 250 615 281
rect 487 247 615 250
rect 512 215 615 247
rect 695 219 729 315
rect 286 17 341 127
rect 512 119 546 215
rect 695 159 754 219
rect 463 53 546 119
rect 591 153 754 159
rect 591 125 729 153
rect 591 61 625 125
rect 674 17 740 89
rect 846 61 891 493
rect 927 450 1093 484
rect 925 315 1025 391
rect 925 141 969 315
rect 1059 281 1093 450
rect 1141 441 1217 527
rect 1277 407 1311 475
rect 1127 357 1397 407
rect 1435 383 1501 527
rect 1710 450 1876 484
rect 1924 451 2000 527
rect 1127 315 1177 357
rect 1279 281 1329 297
rect 1059 247 1329 281
rect 1059 239 1143 247
rect 1005 129 1075 203
rect 1109 93 1143 239
rect 1285 231 1329 247
rect 1363 213 1397 357
rect 1431 283 1632 331
rect 1672 315 1719 397
rect 1431 247 1497 283
rect 1767 261 1808 381
rect 1559 213 1625 247
rect 1177 193 1243 213
rect 1177 187 1259 193
rect 1177 153 1225 187
rect 1363 179 1625 213
rect 1684 225 1808 261
rect 1842 281 1876 450
rect 2048 417 2082 475
rect 2188 451 2482 527
rect 1910 383 2482 417
rect 1910 315 1960 383
rect 1842 247 2112 281
rect 1363 153 1407 179
rect 1177 147 1259 153
rect 1341 119 1407 153
rect 940 53 1143 93
rect 1177 17 1211 105
rect 1245 85 1311 101
rect 1441 85 1475 143
rect 1684 141 1741 225
rect 1842 93 1876 247
rect 2068 215 2112 247
rect 1951 187 2026 213
rect 1951 153 1961 187
rect 1995 153 2026 187
rect 2146 156 2182 383
rect 1951 147 2026 153
rect 2116 119 2182 156
rect 2216 315 2385 349
rect 2216 185 2271 315
rect 2448 265 2482 383
rect 2448 199 2496 265
rect 2216 151 2369 185
rect 1245 51 1475 85
rect 1529 17 1595 93
rect 1723 53 1876 93
rect 1912 17 1964 105
rect 2016 85 2082 109
rect 2216 85 2250 117
rect 2016 51 2250 85
rect 2324 53 2369 151
rect 2416 17 2482 161
rect 2600 299 2647 527
rect 2691 265 2754 483
rect 2790 353 2849 527
rect 2967 299 3015 527
rect 2691 199 2858 265
rect 2600 17 2647 177
rect 2691 51 2754 199
rect 2790 17 2849 109
rect 2967 17 3015 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 1225 153 1259 187
rect 1961 153 1995 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
<< metal1 >>
rect 0 561 3036 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 0 496 3036 527
rect 1213 187 1271 193
rect 1213 153 1225 187
rect 1259 184 1271 187
rect 1949 187 2007 193
rect 1949 184 1961 187
rect 1259 156 1961 184
rect 1259 153 1271 156
rect 1213 147 1271 153
rect 1949 153 1961 156
rect 1995 153 2007 187
rect 1949 147 2007 153
rect 0 17 3036 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
rect 0 -48 3036 -17
<< obsm1 >>
rect 201 388 259 397
rect 937 388 995 397
rect 1673 388 1731 397
rect 201 360 1731 388
rect 201 351 259 360
rect 937 351 995 360
rect 1673 351 1731 360
rect 1581 320 1639 329
rect 2225 320 2283 329
rect 1581 292 2283 320
rect 1581 283 1639 292
rect 2225 283 2283 292
rect 569 252 627 261
rect 845 252 903 261
rect 1673 252 1731 261
rect 569 224 903 252
rect 569 215 627 224
rect 845 215 903 224
rect 1044 224 1731 252
rect 1044 193 1087 224
rect 1673 215 1731 224
rect 109 184 167 193
rect 1029 184 1087 193
rect 109 156 1087 184
rect 109 147 167 156
rect 1029 147 1087 156
<< labels >>
rlabel locali s 17 195 87 325 6 CLK_N
port 1 nsew clock input
rlabel locali s 765 265 805 475 6 D
port 2 nsew signal input
rlabel locali s 2318 219 2414 265 6 RESET_B
port 3 nsew signal input
rlabel locali s 283 205 339 337 6 SCD
port 4 nsew signal input
rlabel locali s 387 69 429 153 6 SCE
port 5 nsew signal input
rlabel locali s 387 153 467 219 6 SCE
port 5 nsew signal input
rlabel locali s 387 219 431 339 6 SCE
port 5 nsew signal input
rlabel metal1 s 1949 147 2007 156 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 147 1271 156 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 156 2007 184 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1949 184 2007 193 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 184 1271 193 6 SET_B
port 6 nsew signal input
rlabel metal1 s 0 -48 3036 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1 21 3035 157 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 2016 157 3035 201 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1241 157 1695 201 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 2398 201 3035 203 6 VNB
port 8 nsew ground bidirectional
rlabel nwell s -38 261 3074 582 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 496 3036 592 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 2883 51 2933 165 6 Q
port 11 nsew signal output
rlabel locali s 2892 165 2933 289 6 Q
port 11 nsew signal output
rlabel locali s 2883 289 2933 493 6 Q
port 11 nsew signal output
rlabel locali s 2516 51 2566 143 6 Q_N
port 12 nsew signal output
rlabel locali s 2532 143 2566 326 6 Q_N
port 12 nsew signal output
rlabel locali s 2516 326 2566 493 6 Q_N
port 12 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3036 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 218634
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 195260
<< end >>
