magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 775 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 247 177
rect 193 127 203 161
rect 237 127 247 161
rect 193 93 247 127
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 93 331 177
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 161 415 177
rect 361 127 371 161
rect 405 127 415 161
rect 361 93 415 127
rect 361 59 371 93
rect 405 59 415 93
rect 361 47 415 59
rect 445 161 499 177
rect 445 127 455 161
rect 489 127 499 161
rect 445 47 499 127
rect 529 93 583 177
rect 529 59 539 93
rect 573 59 583 93
rect 529 47 583 59
rect 613 161 667 177
rect 613 127 623 161
rect 657 127 667 161
rect 613 47 667 127
rect 697 161 749 177
rect 697 127 707 161
rect 741 127 749 161
rect 697 93 749 127
rect 697 59 707 93
rect 741 59 749 93
rect 697 47 749 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 349 499 383
rect 445 315 455 349
rect 489 315 499 349
rect 445 297 499 315
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 349 667 383
rect 613 315 623 349
rect 657 315 667 349
rect 613 297 667 315
rect 697 485 749 497
rect 697 451 707 485
rect 741 451 749 485
rect 697 417 749 451
rect 697 383 707 417
rect 741 383 749 417
rect 697 297 749 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 203 127 237 161
rect 203 59 237 93
rect 287 59 321 93
rect 371 127 405 161
rect 371 59 405 93
rect 455 127 489 161
rect 539 59 573 93
rect 623 127 657 161
rect 707 127 741 161
rect 707 59 741 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 455 451 489 485
rect 455 383 489 417
rect 455 315 489 349
rect 539 451 573 485
rect 539 383 573 417
rect 623 451 657 485
rect 623 383 657 417
rect 623 315 657 349
rect 707 451 741 485
rect 707 383 741 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 22 249 361 265
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 361 249
rect 22 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 415 249 697 265
rect 415 215 539 249
rect 573 215 623 249
rect 657 215 697 249
rect 415 199 697 215
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
<< polycont >>
rect 38 215 72 249
rect 119 215 153 249
rect 203 215 237 249
rect 287 215 321 249
rect 539 215 573 249
rect 623 215 657 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 405 527
rect 371 417 405 451
rect 371 367 405 383
rect 439 485 505 493
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 439 349 505 383
rect 539 485 573 527
rect 539 417 573 451
rect 539 367 573 383
rect 607 485 673 493
rect 607 451 623 485
rect 657 451 673 485
rect 607 417 673 451
rect 607 383 623 417
rect 657 383 673 417
rect 439 333 455 349
rect 321 315 455 333
rect 489 333 505 349
rect 607 349 673 383
rect 707 485 757 527
rect 741 451 757 485
rect 707 417 757 451
rect 741 383 757 417
rect 707 367 757 383
rect 607 333 623 349
rect 489 315 623 333
rect 657 315 673 349
rect 103 299 673 315
rect 22 249 346 265
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 346 249
rect 382 215 489 299
rect 523 249 811 265
rect 523 215 539 249
rect 573 215 623 249
rect 657 215 811 249
rect 18 161 405 181
rect 18 127 35 161
rect 69 143 203 161
rect 69 127 85 143
rect 18 93 85 127
rect 187 127 203 143
rect 237 143 371 161
rect 237 127 253 143
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 119 93 153 109
rect 119 17 153 59
rect 187 93 253 127
rect 355 127 371 143
rect 439 161 489 215
rect 707 161 757 177
rect 439 127 455 161
rect 489 127 623 161
rect 657 127 673 161
rect 741 127 757 161
rect 187 59 203 93
rect 237 59 253 93
rect 187 51 253 59
rect 287 93 321 109
rect 287 17 321 59
rect 355 93 405 127
rect 707 93 757 127
rect 355 59 371 93
rect 405 59 539 93
rect 573 59 707 93
rect 741 59 757 93
rect 355 51 757 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 398 289 432 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 674 221 708 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand2_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1717208
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1709626
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
