magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< poly >>
rect 1671 435 1701 896
rect 2295 559 2325 896
rect 2919 683 2949 896
rect 3543 807 3573 896
rect 3525 791 3591 807
rect 3525 757 3541 791
rect 3575 757 3591 791
rect 3525 741 3591 757
rect 2901 667 2967 683
rect 2901 633 2917 667
rect 2951 633 2967 667
rect 2901 617 2967 633
rect 2277 543 2343 559
rect 2277 509 2293 543
rect 2327 509 2343 543
rect 2277 493 2343 509
rect 4167 435 4197 896
rect 4791 559 4821 896
rect 5415 683 5445 896
rect 6039 807 6069 896
rect 6021 791 6087 807
rect 6021 757 6037 791
rect 6071 757 6087 791
rect 6021 741 6087 757
rect 5397 667 5463 683
rect 5397 633 5413 667
rect 5447 633 5463 667
rect 5397 617 5463 633
rect 4773 543 4839 559
rect 4773 509 4789 543
rect 4823 509 4839 543
rect 4773 493 4839 509
rect 6663 435 6693 896
rect 7287 559 7317 896
rect 7911 683 7941 896
rect 8535 807 8565 896
rect 8517 791 8583 807
rect 8517 757 8533 791
rect 8567 757 8583 791
rect 8517 741 8583 757
rect 7893 667 7959 683
rect 7893 633 7909 667
rect 7943 633 7959 667
rect 7893 617 7959 633
rect 7269 543 7335 559
rect 7269 509 7285 543
rect 7319 509 7335 543
rect 7269 493 7335 509
rect 9159 435 9189 896
rect 9783 559 9813 896
rect 10407 683 10437 896
rect 11031 807 11061 896
rect 11013 791 11079 807
rect 11013 757 11029 791
rect 11063 757 11079 791
rect 11013 741 11079 757
rect 10389 667 10455 683
rect 10389 633 10405 667
rect 10439 633 10455 667
rect 10389 617 10455 633
rect 9765 543 9831 559
rect 9765 509 9781 543
rect 9815 509 9831 543
rect 9765 493 9831 509
rect 11655 435 11685 896
rect 12279 559 12309 896
rect 12903 683 12933 896
rect 13527 807 13557 896
rect 13509 791 13575 807
rect 13509 757 13525 791
rect 13559 757 13575 791
rect 13509 741 13575 757
rect 12885 667 12951 683
rect 12885 633 12901 667
rect 12935 633 12951 667
rect 12885 617 12951 633
rect 12261 543 12327 559
rect 12261 509 12277 543
rect 12311 509 12327 543
rect 12261 493 12327 509
rect 14151 435 14181 896
rect 14775 559 14805 896
rect 15399 683 15429 896
rect 16023 807 16053 896
rect 16005 791 16071 807
rect 16005 757 16021 791
rect 16055 757 16071 791
rect 16005 741 16071 757
rect 15381 667 15447 683
rect 15381 633 15397 667
rect 15431 633 15447 667
rect 15381 617 15447 633
rect 14757 543 14823 559
rect 14757 509 14773 543
rect 14807 509 14823 543
rect 14757 493 14823 509
rect 16647 435 16677 896
rect 17271 559 17301 896
rect 17895 683 17925 896
rect 18519 807 18549 896
rect 18501 791 18567 807
rect 18501 757 18517 791
rect 18551 757 18567 791
rect 18501 741 18567 757
rect 17877 667 17943 683
rect 17877 633 17893 667
rect 17927 633 17943 667
rect 17877 617 17943 633
rect 17253 543 17319 559
rect 17253 509 17269 543
rect 17303 509 17319 543
rect 17253 493 17319 509
rect 19143 435 19173 896
rect 19767 559 19797 896
rect 20391 683 20421 896
rect 21015 807 21045 896
rect 20997 791 21063 807
rect 20997 757 21013 791
rect 21047 757 21063 791
rect 20997 741 21063 757
rect 20373 667 20439 683
rect 20373 633 20389 667
rect 20423 633 20439 667
rect 20373 617 20439 633
rect 19749 543 19815 559
rect 19749 509 19765 543
rect 19799 509 19815 543
rect 19749 493 19815 509
rect 21639 435 21669 896
rect 22263 559 22293 896
rect 22887 683 22917 896
rect 23511 807 23541 896
rect 23493 791 23559 807
rect 23493 757 23509 791
rect 23543 757 23559 791
rect 23493 741 23559 757
rect 22869 667 22935 683
rect 22869 633 22885 667
rect 22919 633 22935 667
rect 22869 617 22935 633
rect 22245 543 22311 559
rect 22245 509 22261 543
rect 22295 509 22311 543
rect 22245 493 22311 509
rect 24135 435 24165 896
rect 24759 559 24789 896
rect 25383 683 25413 896
rect 26007 807 26037 896
rect 25989 791 26055 807
rect 25989 757 26005 791
rect 26039 757 26055 791
rect 25989 741 26055 757
rect 25365 667 25431 683
rect 25365 633 25381 667
rect 25415 633 25431 667
rect 25365 617 25431 633
rect 24741 543 24807 559
rect 24741 509 24757 543
rect 24791 509 24807 543
rect 24741 493 24807 509
rect 26631 435 26661 896
rect 27255 559 27285 896
rect 27879 683 27909 896
rect 28503 807 28533 896
rect 28485 791 28551 807
rect 28485 757 28501 791
rect 28535 757 28551 791
rect 28485 741 28551 757
rect 27861 667 27927 683
rect 27861 633 27877 667
rect 27911 633 27927 667
rect 27861 617 27927 633
rect 27237 543 27303 559
rect 27237 509 27253 543
rect 27287 509 27303 543
rect 27237 493 27303 509
rect 29127 435 29157 896
rect 29751 559 29781 896
rect 30375 683 30405 896
rect 30999 807 31029 896
rect 30981 791 31047 807
rect 30981 757 30997 791
rect 31031 757 31047 791
rect 30981 741 31047 757
rect 30357 667 30423 683
rect 30357 633 30373 667
rect 30407 633 30423 667
rect 30357 617 30423 633
rect 29733 543 29799 559
rect 29733 509 29749 543
rect 29783 509 29799 543
rect 29733 493 29799 509
rect 31623 435 31653 896
rect 32247 559 32277 896
rect 32871 683 32901 896
rect 33495 807 33525 896
rect 33477 791 33543 807
rect 33477 757 33493 791
rect 33527 757 33543 791
rect 33477 741 33543 757
rect 32853 667 32919 683
rect 32853 633 32869 667
rect 32903 633 32919 667
rect 32853 617 32919 633
rect 32229 543 32295 559
rect 32229 509 32245 543
rect 32279 509 32295 543
rect 32229 493 32295 509
rect 34119 435 34149 896
rect 34743 559 34773 896
rect 35367 683 35397 896
rect 35991 807 36021 896
rect 35973 791 36039 807
rect 35973 757 35989 791
rect 36023 757 36039 791
rect 35973 741 36039 757
rect 35349 667 35415 683
rect 35349 633 35365 667
rect 35399 633 35415 667
rect 35349 617 35415 633
rect 34725 543 34791 559
rect 34725 509 34741 543
rect 34775 509 34791 543
rect 34725 493 34791 509
rect 36615 435 36645 896
rect 37239 559 37269 896
rect 37863 683 37893 896
rect 38487 807 38517 896
rect 38469 791 38535 807
rect 38469 757 38485 791
rect 38519 757 38535 791
rect 38469 741 38535 757
rect 37845 667 37911 683
rect 37845 633 37861 667
rect 37895 633 37911 667
rect 37845 617 37911 633
rect 37221 543 37287 559
rect 37221 509 37237 543
rect 37271 509 37287 543
rect 37221 493 37287 509
rect 39111 435 39141 896
rect 39735 559 39765 896
rect 40359 683 40389 896
rect 40983 807 41013 896
rect 40965 791 41031 807
rect 40965 757 40981 791
rect 41015 757 41031 791
rect 40965 741 41031 757
rect 40341 667 40407 683
rect 40341 633 40357 667
rect 40391 633 40407 667
rect 40341 617 40407 633
rect 39717 543 39783 559
rect 39717 509 39733 543
rect 39767 509 39783 543
rect 39717 493 39783 509
rect 41607 435 41637 896
rect 42231 559 42261 896
rect 42855 683 42885 896
rect 43479 807 43509 896
rect 43461 791 43527 807
rect 43461 757 43477 791
rect 43511 757 43527 791
rect 43461 741 43527 757
rect 42837 667 42903 683
rect 42837 633 42853 667
rect 42887 633 42903 667
rect 42837 617 42903 633
rect 42213 543 42279 559
rect 42213 509 42229 543
rect 42263 509 42279 543
rect 42213 493 42279 509
rect 44103 435 44133 896
rect 44727 559 44757 896
rect 45351 683 45381 896
rect 45975 807 46005 896
rect 45957 791 46023 807
rect 45957 757 45973 791
rect 46007 757 46023 791
rect 45957 741 46023 757
rect 45333 667 45399 683
rect 45333 633 45349 667
rect 45383 633 45399 667
rect 45333 617 45399 633
rect 44709 543 44775 559
rect 44709 509 44725 543
rect 44759 509 44775 543
rect 44709 493 44775 509
rect 46599 435 46629 896
rect 47223 559 47253 896
rect 47847 683 47877 896
rect 48471 807 48501 896
rect 48453 791 48519 807
rect 48453 757 48469 791
rect 48503 757 48519 791
rect 48453 741 48519 757
rect 47829 667 47895 683
rect 47829 633 47845 667
rect 47879 633 47895 667
rect 47829 617 47895 633
rect 47205 543 47271 559
rect 47205 509 47221 543
rect 47255 509 47271 543
rect 47205 493 47271 509
rect 49095 435 49125 896
rect 49719 559 49749 896
rect 50343 683 50373 896
rect 50967 807 50997 896
rect 50949 791 51015 807
rect 50949 757 50965 791
rect 50999 757 51015 791
rect 50949 741 51015 757
rect 50325 667 50391 683
rect 50325 633 50341 667
rect 50375 633 50391 667
rect 50325 617 50391 633
rect 49701 543 49767 559
rect 49701 509 49717 543
rect 49751 509 49767 543
rect 49701 493 49767 509
rect 51591 435 51621 896
rect 52215 559 52245 896
rect 52839 683 52869 896
rect 53463 807 53493 896
rect 53445 791 53511 807
rect 53445 757 53461 791
rect 53495 757 53511 791
rect 53445 741 53511 757
rect 52821 667 52887 683
rect 52821 633 52837 667
rect 52871 633 52887 667
rect 52821 617 52887 633
rect 52197 543 52263 559
rect 52197 509 52213 543
rect 52247 509 52263 543
rect 52197 493 52263 509
rect 54087 435 54117 896
rect 54711 559 54741 896
rect 55335 683 55365 896
rect 55959 807 55989 896
rect 55941 791 56007 807
rect 55941 757 55957 791
rect 55991 757 56007 791
rect 55941 741 56007 757
rect 55317 667 55383 683
rect 55317 633 55333 667
rect 55367 633 55383 667
rect 55317 617 55383 633
rect 54693 543 54759 559
rect 54693 509 54709 543
rect 54743 509 54759 543
rect 54693 493 54759 509
rect 56583 435 56613 896
rect 57207 559 57237 896
rect 57831 683 57861 896
rect 58455 807 58485 896
rect 58437 791 58503 807
rect 58437 757 58453 791
rect 58487 757 58503 791
rect 58437 741 58503 757
rect 57813 667 57879 683
rect 57813 633 57829 667
rect 57863 633 57879 667
rect 57813 617 57879 633
rect 57189 543 57255 559
rect 57189 509 57205 543
rect 57239 509 57255 543
rect 57189 493 57255 509
rect 59079 435 59109 896
rect 59703 559 59733 896
rect 60327 683 60357 896
rect 60951 807 60981 896
rect 60933 791 60999 807
rect 60933 757 60949 791
rect 60983 757 60999 791
rect 60933 741 60999 757
rect 60309 667 60375 683
rect 60309 633 60325 667
rect 60359 633 60375 667
rect 60309 617 60375 633
rect 59685 543 59751 559
rect 59685 509 59701 543
rect 59735 509 59751 543
rect 59685 493 59751 509
rect 61575 435 61605 896
rect 62199 559 62229 896
rect 62823 683 62853 896
rect 63447 807 63477 896
rect 63429 791 63495 807
rect 63429 757 63445 791
rect 63479 757 63495 791
rect 63429 741 63495 757
rect 62805 667 62871 683
rect 62805 633 62821 667
rect 62855 633 62871 667
rect 62805 617 62871 633
rect 62181 543 62247 559
rect 62181 509 62197 543
rect 62231 509 62247 543
rect 62181 493 62247 509
rect 64071 435 64101 896
rect 64695 559 64725 896
rect 65319 683 65349 896
rect 65943 807 65973 896
rect 65925 791 65991 807
rect 65925 757 65941 791
rect 65975 757 65991 791
rect 65925 741 65991 757
rect 65301 667 65367 683
rect 65301 633 65317 667
rect 65351 633 65367 667
rect 65301 617 65367 633
rect 64677 543 64743 559
rect 64677 509 64693 543
rect 64727 509 64743 543
rect 64677 493 64743 509
rect 66567 435 66597 896
rect 67191 559 67221 896
rect 67815 683 67845 896
rect 68439 807 68469 896
rect 68421 791 68487 807
rect 68421 757 68437 791
rect 68471 757 68487 791
rect 68421 741 68487 757
rect 67797 667 67863 683
rect 67797 633 67813 667
rect 67847 633 67863 667
rect 67797 617 67863 633
rect 67173 543 67239 559
rect 67173 509 67189 543
rect 67223 509 67239 543
rect 67173 493 67239 509
rect 69063 435 69093 896
rect 69687 559 69717 896
rect 70311 683 70341 896
rect 70935 807 70965 896
rect 70917 791 70983 807
rect 70917 757 70933 791
rect 70967 757 70983 791
rect 70917 741 70983 757
rect 70293 667 70359 683
rect 70293 633 70309 667
rect 70343 633 70359 667
rect 70293 617 70359 633
rect 69669 543 69735 559
rect 69669 509 69685 543
rect 69719 509 69735 543
rect 69669 493 69735 509
rect 71559 435 71589 896
rect 72183 559 72213 896
rect 72807 683 72837 896
rect 73431 807 73461 896
rect 73413 791 73479 807
rect 73413 757 73429 791
rect 73463 757 73479 791
rect 73413 741 73479 757
rect 72789 667 72855 683
rect 72789 633 72805 667
rect 72839 633 72855 667
rect 72789 617 72855 633
rect 72165 543 72231 559
rect 72165 509 72181 543
rect 72215 509 72231 543
rect 72165 493 72231 509
rect 74055 435 74085 896
rect 74679 559 74709 896
rect 75303 683 75333 896
rect 75927 807 75957 896
rect 75909 791 75975 807
rect 75909 757 75925 791
rect 75959 757 75975 791
rect 75909 741 75975 757
rect 75285 667 75351 683
rect 75285 633 75301 667
rect 75335 633 75351 667
rect 75285 617 75351 633
rect 74661 543 74727 559
rect 74661 509 74677 543
rect 74711 509 74727 543
rect 74661 493 74727 509
rect 76551 435 76581 896
rect 77175 559 77205 896
rect 77799 683 77829 896
rect 78423 807 78453 896
rect 78405 791 78471 807
rect 78405 757 78421 791
rect 78455 757 78471 791
rect 78405 741 78471 757
rect 77781 667 77847 683
rect 77781 633 77797 667
rect 77831 633 77847 667
rect 77781 617 77847 633
rect 77157 543 77223 559
rect 77157 509 77173 543
rect 77207 509 77223 543
rect 77157 493 77223 509
rect 79047 435 79077 896
rect 79671 559 79701 896
rect 80295 683 80325 896
rect 80919 807 80949 896
rect 80901 791 80967 807
rect 80901 757 80917 791
rect 80951 757 80967 791
rect 80901 741 80967 757
rect 80277 667 80343 683
rect 80277 633 80293 667
rect 80327 633 80343 667
rect 80277 617 80343 633
rect 79653 543 79719 559
rect 79653 509 79669 543
rect 79703 509 79719 543
rect 79653 493 79719 509
rect 1653 419 1719 435
rect 1653 385 1669 419
rect 1703 385 1719 419
rect 1653 369 1719 385
rect 4149 419 4215 435
rect 4149 385 4165 419
rect 4199 385 4215 419
rect 4149 369 4215 385
rect 6645 419 6711 435
rect 6645 385 6661 419
rect 6695 385 6711 419
rect 6645 369 6711 385
rect 9141 419 9207 435
rect 9141 385 9157 419
rect 9191 385 9207 419
rect 9141 369 9207 385
rect 11637 419 11703 435
rect 11637 385 11653 419
rect 11687 385 11703 419
rect 11637 369 11703 385
rect 14133 419 14199 435
rect 14133 385 14149 419
rect 14183 385 14199 419
rect 14133 369 14199 385
rect 16629 419 16695 435
rect 16629 385 16645 419
rect 16679 385 16695 419
rect 16629 369 16695 385
rect 19125 419 19191 435
rect 19125 385 19141 419
rect 19175 385 19191 419
rect 19125 369 19191 385
rect 21621 419 21687 435
rect 21621 385 21637 419
rect 21671 385 21687 419
rect 21621 369 21687 385
rect 24117 419 24183 435
rect 24117 385 24133 419
rect 24167 385 24183 419
rect 24117 369 24183 385
rect 26613 419 26679 435
rect 26613 385 26629 419
rect 26663 385 26679 419
rect 26613 369 26679 385
rect 29109 419 29175 435
rect 29109 385 29125 419
rect 29159 385 29175 419
rect 29109 369 29175 385
rect 31605 419 31671 435
rect 31605 385 31621 419
rect 31655 385 31671 419
rect 31605 369 31671 385
rect 34101 419 34167 435
rect 34101 385 34117 419
rect 34151 385 34167 419
rect 34101 369 34167 385
rect 36597 419 36663 435
rect 36597 385 36613 419
rect 36647 385 36663 419
rect 36597 369 36663 385
rect 39093 419 39159 435
rect 39093 385 39109 419
rect 39143 385 39159 419
rect 39093 369 39159 385
rect 41589 419 41655 435
rect 41589 385 41605 419
rect 41639 385 41655 419
rect 41589 369 41655 385
rect 44085 419 44151 435
rect 44085 385 44101 419
rect 44135 385 44151 419
rect 44085 369 44151 385
rect 46581 419 46647 435
rect 46581 385 46597 419
rect 46631 385 46647 419
rect 46581 369 46647 385
rect 49077 419 49143 435
rect 49077 385 49093 419
rect 49127 385 49143 419
rect 49077 369 49143 385
rect 51573 419 51639 435
rect 51573 385 51589 419
rect 51623 385 51639 419
rect 51573 369 51639 385
rect 54069 419 54135 435
rect 54069 385 54085 419
rect 54119 385 54135 419
rect 54069 369 54135 385
rect 56565 419 56631 435
rect 56565 385 56581 419
rect 56615 385 56631 419
rect 56565 369 56631 385
rect 59061 419 59127 435
rect 59061 385 59077 419
rect 59111 385 59127 419
rect 59061 369 59127 385
rect 61557 419 61623 435
rect 61557 385 61573 419
rect 61607 385 61623 419
rect 61557 369 61623 385
rect 64053 419 64119 435
rect 64053 385 64069 419
rect 64103 385 64119 419
rect 64053 369 64119 385
rect 66549 419 66615 435
rect 66549 385 66565 419
rect 66599 385 66615 419
rect 66549 369 66615 385
rect 69045 419 69111 435
rect 69045 385 69061 419
rect 69095 385 69111 419
rect 69045 369 69111 385
rect 71541 419 71607 435
rect 71541 385 71557 419
rect 71591 385 71607 419
rect 71541 369 71607 385
rect 74037 419 74103 435
rect 74037 385 74053 419
rect 74087 385 74103 419
rect 74037 369 74103 385
rect 76533 419 76599 435
rect 76533 385 76549 419
rect 76583 385 76599 419
rect 76533 369 76599 385
rect 79029 419 79095 435
rect 79029 385 79045 419
rect 79079 385 79095 419
rect 79029 369 79095 385
<< polycont >>
rect 3541 757 3575 791
rect 2917 633 2951 667
rect 2293 509 2327 543
rect 6037 757 6071 791
rect 5413 633 5447 667
rect 4789 509 4823 543
rect 8533 757 8567 791
rect 7909 633 7943 667
rect 7285 509 7319 543
rect 11029 757 11063 791
rect 10405 633 10439 667
rect 9781 509 9815 543
rect 13525 757 13559 791
rect 12901 633 12935 667
rect 12277 509 12311 543
rect 16021 757 16055 791
rect 15397 633 15431 667
rect 14773 509 14807 543
rect 18517 757 18551 791
rect 17893 633 17927 667
rect 17269 509 17303 543
rect 21013 757 21047 791
rect 20389 633 20423 667
rect 19765 509 19799 543
rect 23509 757 23543 791
rect 22885 633 22919 667
rect 22261 509 22295 543
rect 26005 757 26039 791
rect 25381 633 25415 667
rect 24757 509 24791 543
rect 28501 757 28535 791
rect 27877 633 27911 667
rect 27253 509 27287 543
rect 30997 757 31031 791
rect 30373 633 30407 667
rect 29749 509 29783 543
rect 33493 757 33527 791
rect 32869 633 32903 667
rect 32245 509 32279 543
rect 35989 757 36023 791
rect 35365 633 35399 667
rect 34741 509 34775 543
rect 38485 757 38519 791
rect 37861 633 37895 667
rect 37237 509 37271 543
rect 40981 757 41015 791
rect 40357 633 40391 667
rect 39733 509 39767 543
rect 43477 757 43511 791
rect 42853 633 42887 667
rect 42229 509 42263 543
rect 45973 757 46007 791
rect 45349 633 45383 667
rect 44725 509 44759 543
rect 48469 757 48503 791
rect 47845 633 47879 667
rect 47221 509 47255 543
rect 50965 757 50999 791
rect 50341 633 50375 667
rect 49717 509 49751 543
rect 53461 757 53495 791
rect 52837 633 52871 667
rect 52213 509 52247 543
rect 55957 757 55991 791
rect 55333 633 55367 667
rect 54709 509 54743 543
rect 58453 757 58487 791
rect 57829 633 57863 667
rect 57205 509 57239 543
rect 60949 757 60983 791
rect 60325 633 60359 667
rect 59701 509 59735 543
rect 63445 757 63479 791
rect 62821 633 62855 667
rect 62197 509 62231 543
rect 65941 757 65975 791
rect 65317 633 65351 667
rect 64693 509 64727 543
rect 68437 757 68471 791
rect 67813 633 67847 667
rect 67189 509 67223 543
rect 70933 757 70967 791
rect 70309 633 70343 667
rect 69685 509 69719 543
rect 73429 757 73463 791
rect 72805 633 72839 667
rect 72181 509 72215 543
rect 75925 757 75959 791
rect 75301 633 75335 667
rect 74677 509 74711 543
rect 78421 757 78455 791
rect 77797 633 77831 667
rect 77173 509 77207 543
rect 80917 757 80951 791
rect 80293 633 80327 667
rect 79669 509 79703 543
rect 1669 385 1703 419
rect 4165 385 4199 419
rect 6661 385 6695 419
rect 9157 385 9191 419
rect 11653 385 11687 419
rect 14149 385 14183 419
rect 16645 385 16679 419
rect 19141 385 19175 419
rect 21637 385 21671 419
rect 24133 385 24167 419
rect 26629 385 26663 419
rect 29125 385 29159 419
rect 31621 385 31655 419
rect 34117 385 34151 419
rect 36613 385 36647 419
rect 39109 385 39143 419
rect 41605 385 41639 419
rect 44101 385 44135 419
rect 46597 385 46631 419
rect 49093 385 49127 419
rect 51589 385 51623 419
rect 54085 385 54119 419
rect 56581 385 56615 419
rect 59077 385 59111 419
rect 61573 385 61607 419
rect 64069 385 64103 419
rect 66565 385 66599 419
rect 69061 385 69095 419
rect 71557 385 71591 419
rect 74053 385 74087 419
rect 76549 385 76583 419
rect 79045 385 79079 419
<< locali >>
rect 3541 791 3575 807
rect 3541 741 3575 757
rect 6037 791 6071 807
rect 6037 741 6071 757
rect 8533 791 8567 807
rect 8533 741 8567 757
rect 11029 791 11063 807
rect 11029 741 11063 757
rect 13525 791 13559 807
rect 13525 741 13559 757
rect 16021 791 16055 807
rect 16021 741 16055 757
rect 18517 791 18551 807
rect 18517 741 18551 757
rect 21013 791 21047 807
rect 21013 741 21047 757
rect 23509 791 23543 807
rect 23509 741 23543 757
rect 26005 791 26039 807
rect 26005 741 26039 757
rect 28501 791 28535 807
rect 28501 741 28535 757
rect 30997 791 31031 807
rect 30997 741 31031 757
rect 33493 791 33527 807
rect 33493 741 33527 757
rect 35989 791 36023 807
rect 35989 741 36023 757
rect 38485 791 38519 807
rect 38485 741 38519 757
rect 40981 791 41015 807
rect 40981 741 41015 757
rect 43477 791 43511 807
rect 43477 741 43511 757
rect 45973 791 46007 807
rect 45973 741 46007 757
rect 48469 791 48503 807
rect 48469 741 48503 757
rect 50965 791 50999 807
rect 50965 741 50999 757
rect 53461 791 53495 807
rect 53461 741 53495 757
rect 55957 791 55991 807
rect 55957 741 55991 757
rect 58453 791 58487 807
rect 58453 741 58487 757
rect 60949 791 60983 807
rect 60949 741 60983 757
rect 63445 791 63479 807
rect 63445 741 63479 757
rect 65941 791 65975 807
rect 65941 741 65975 757
rect 68437 791 68471 807
rect 68437 741 68471 757
rect 70933 791 70967 807
rect 70933 741 70967 757
rect 73429 791 73463 807
rect 73429 741 73463 757
rect 75925 791 75959 807
rect 75925 741 75959 757
rect 78421 791 78455 807
rect 78421 741 78455 757
rect 80917 791 80951 807
rect 80917 741 80951 757
rect 2917 667 2951 683
rect 2917 617 2951 633
rect 5413 667 5447 683
rect 5413 617 5447 633
rect 7909 667 7943 683
rect 7909 617 7943 633
rect 10405 667 10439 683
rect 10405 617 10439 633
rect 12901 667 12935 683
rect 12901 617 12935 633
rect 15397 667 15431 683
rect 15397 617 15431 633
rect 17893 667 17927 683
rect 17893 617 17927 633
rect 20389 667 20423 683
rect 20389 617 20423 633
rect 22885 667 22919 683
rect 22885 617 22919 633
rect 25381 667 25415 683
rect 25381 617 25415 633
rect 27877 667 27911 683
rect 27877 617 27911 633
rect 30373 667 30407 683
rect 30373 617 30407 633
rect 32869 667 32903 683
rect 32869 617 32903 633
rect 35365 667 35399 683
rect 35365 617 35399 633
rect 37861 667 37895 683
rect 37861 617 37895 633
rect 40357 667 40391 683
rect 40357 617 40391 633
rect 42853 667 42887 683
rect 42853 617 42887 633
rect 45349 667 45383 683
rect 45349 617 45383 633
rect 47845 667 47879 683
rect 47845 617 47879 633
rect 50341 667 50375 683
rect 50341 617 50375 633
rect 52837 667 52871 683
rect 52837 617 52871 633
rect 55333 667 55367 683
rect 55333 617 55367 633
rect 57829 667 57863 683
rect 57829 617 57863 633
rect 60325 667 60359 683
rect 60325 617 60359 633
rect 62821 667 62855 683
rect 62821 617 62855 633
rect 65317 667 65351 683
rect 65317 617 65351 633
rect 67813 667 67847 683
rect 67813 617 67847 633
rect 70309 667 70343 683
rect 70309 617 70343 633
rect 72805 667 72839 683
rect 72805 617 72839 633
rect 75301 667 75335 683
rect 75301 617 75335 633
rect 77797 667 77831 683
rect 77797 617 77831 633
rect 80293 667 80327 683
rect 80293 617 80327 633
rect 2293 543 2327 559
rect 2293 493 2327 509
rect 4789 543 4823 559
rect 4789 493 4823 509
rect 7285 543 7319 559
rect 7285 493 7319 509
rect 9781 543 9815 559
rect 9781 493 9815 509
rect 12277 543 12311 559
rect 12277 493 12311 509
rect 14773 543 14807 559
rect 14773 493 14807 509
rect 17269 543 17303 559
rect 17269 493 17303 509
rect 19765 543 19799 559
rect 19765 493 19799 509
rect 22261 543 22295 559
rect 22261 493 22295 509
rect 24757 543 24791 559
rect 24757 493 24791 509
rect 27253 543 27287 559
rect 27253 493 27287 509
rect 29749 543 29783 559
rect 29749 493 29783 509
rect 32245 543 32279 559
rect 32245 493 32279 509
rect 34741 543 34775 559
rect 34741 493 34775 509
rect 37237 543 37271 559
rect 37237 493 37271 509
rect 39733 543 39767 559
rect 39733 493 39767 509
rect 42229 543 42263 559
rect 42229 493 42263 509
rect 44725 543 44759 559
rect 44725 493 44759 509
rect 47221 543 47255 559
rect 47221 493 47255 509
rect 49717 543 49751 559
rect 49717 493 49751 509
rect 52213 543 52247 559
rect 52213 493 52247 509
rect 54709 543 54743 559
rect 54709 493 54743 509
rect 57205 543 57239 559
rect 57205 493 57239 509
rect 59701 543 59735 559
rect 59701 493 59735 509
rect 62197 543 62231 559
rect 62197 493 62231 509
rect 64693 543 64727 559
rect 64693 493 64727 509
rect 67189 543 67223 559
rect 67189 493 67223 509
rect 69685 543 69719 559
rect 69685 493 69719 509
rect 72181 543 72215 559
rect 72181 493 72215 509
rect 74677 543 74711 559
rect 74677 493 74711 509
rect 77173 543 77207 559
rect 77173 493 77207 509
rect 79669 543 79703 559
rect 79669 493 79703 509
rect 1669 419 1703 435
rect 1669 369 1703 385
rect 4165 419 4199 435
rect 4165 369 4199 385
rect 6661 419 6695 435
rect 6661 369 6695 385
rect 9157 419 9191 435
rect 9157 369 9191 385
rect 11653 419 11687 435
rect 11653 369 11687 385
rect 14149 419 14183 435
rect 14149 369 14183 385
rect 16645 419 16679 435
rect 16645 369 16679 385
rect 19141 419 19175 435
rect 19141 369 19175 385
rect 21637 419 21671 435
rect 21637 369 21671 385
rect 24133 419 24167 435
rect 24133 369 24167 385
rect 26629 419 26663 435
rect 26629 369 26663 385
rect 29125 419 29159 435
rect 29125 369 29159 385
rect 31621 419 31655 435
rect 31621 369 31655 385
rect 34117 419 34151 435
rect 34117 369 34151 385
rect 36613 419 36647 435
rect 36613 369 36647 385
rect 39109 419 39143 435
rect 39109 369 39143 385
rect 41605 419 41639 435
rect 41605 369 41639 385
rect 44101 419 44135 435
rect 44101 369 44135 385
rect 46597 419 46631 435
rect 46597 369 46631 385
rect 49093 419 49127 435
rect 49093 369 49127 385
rect 51589 419 51623 435
rect 51589 369 51623 385
rect 54085 419 54119 435
rect 54085 369 54119 385
rect 56581 419 56615 435
rect 56581 369 56615 385
rect 59077 419 59111 435
rect 59077 369 59111 385
rect 61573 419 61607 435
rect 61573 369 61607 385
rect 64069 419 64103 435
rect 64069 369 64103 385
rect 66565 419 66599 435
rect 66565 369 66599 385
rect 69061 419 69095 435
rect 69061 369 69095 385
rect 71557 419 71591 435
rect 71557 369 71591 385
rect 74053 419 74087 435
rect 74053 369 74087 385
rect 76549 419 76583 435
rect 76549 369 76583 385
rect 79045 419 79079 435
rect 79045 369 79079 385
<< viali >>
rect 3541 757 3575 791
rect 6037 757 6071 791
rect 8533 757 8567 791
rect 11029 757 11063 791
rect 13525 757 13559 791
rect 16021 757 16055 791
rect 18517 757 18551 791
rect 21013 757 21047 791
rect 23509 757 23543 791
rect 26005 757 26039 791
rect 28501 757 28535 791
rect 30997 757 31031 791
rect 33493 757 33527 791
rect 35989 757 36023 791
rect 38485 757 38519 791
rect 40981 757 41015 791
rect 43477 757 43511 791
rect 45973 757 46007 791
rect 48469 757 48503 791
rect 50965 757 50999 791
rect 53461 757 53495 791
rect 55957 757 55991 791
rect 58453 757 58487 791
rect 60949 757 60983 791
rect 63445 757 63479 791
rect 65941 757 65975 791
rect 68437 757 68471 791
rect 70933 757 70967 791
rect 73429 757 73463 791
rect 75925 757 75959 791
rect 78421 757 78455 791
rect 80917 757 80951 791
rect 2917 633 2951 667
rect 5413 633 5447 667
rect 7909 633 7943 667
rect 10405 633 10439 667
rect 12901 633 12935 667
rect 15397 633 15431 667
rect 17893 633 17927 667
rect 20389 633 20423 667
rect 22885 633 22919 667
rect 25381 633 25415 667
rect 27877 633 27911 667
rect 30373 633 30407 667
rect 32869 633 32903 667
rect 35365 633 35399 667
rect 37861 633 37895 667
rect 40357 633 40391 667
rect 42853 633 42887 667
rect 45349 633 45383 667
rect 47845 633 47879 667
rect 50341 633 50375 667
rect 52837 633 52871 667
rect 55333 633 55367 667
rect 57829 633 57863 667
rect 60325 633 60359 667
rect 62821 633 62855 667
rect 65317 633 65351 667
rect 67813 633 67847 667
rect 70309 633 70343 667
rect 72805 633 72839 667
rect 75301 633 75335 667
rect 77797 633 77831 667
rect 80293 633 80327 667
rect 2293 509 2327 543
rect 4789 509 4823 543
rect 7285 509 7319 543
rect 9781 509 9815 543
rect 12277 509 12311 543
rect 14773 509 14807 543
rect 17269 509 17303 543
rect 19765 509 19799 543
rect 22261 509 22295 543
rect 24757 509 24791 543
rect 27253 509 27287 543
rect 29749 509 29783 543
rect 32245 509 32279 543
rect 34741 509 34775 543
rect 37237 509 37271 543
rect 39733 509 39767 543
rect 42229 509 42263 543
rect 44725 509 44759 543
rect 47221 509 47255 543
rect 49717 509 49751 543
rect 52213 509 52247 543
rect 54709 509 54743 543
rect 57205 509 57239 543
rect 59701 509 59735 543
rect 62197 509 62231 543
rect 64693 509 64727 543
rect 67189 509 67223 543
rect 69685 509 69719 543
rect 72181 509 72215 543
rect 74677 509 74711 543
rect 77173 509 77207 543
rect 79669 509 79703 543
rect 1669 385 1703 419
rect 4165 385 4199 419
rect 6661 385 6695 419
rect 9157 385 9191 419
rect 11653 385 11687 419
rect 14149 385 14183 419
rect 16645 385 16679 419
rect 19141 385 19175 419
rect 21637 385 21671 419
rect 24133 385 24167 419
rect 26629 385 26663 419
rect 29125 385 29159 419
rect 31621 385 31655 419
rect 34117 385 34151 419
rect 36613 385 36647 419
rect 39109 385 39143 419
rect 41605 385 41639 419
rect 44101 385 44135 419
rect 46597 385 46631 419
rect 49093 385 49127 419
rect 51589 385 51623 419
rect 54085 385 54119 419
rect 56581 385 56615 419
rect 59077 385 59111 419
rect 61573 385 61607 419
rect 64069 385 64103 419
rect 66565 385 66599 419
rect 69061 385 69095 419
rect 71557 385 71591 419
rect 74053 385 74087 419
rect 76549 385 76583 419
rect 79045 385 79079 419
<< metal1 >>
rect 1454 2128 1482 2184
rect 1918 2128 1946 2184
rect 2050 2128 2078 2184
rect 2514 2128 2542 2184
rect 2702 2128 2730 2184
rect 3166 2128 3194 2184
rect 3298 2128 3326 2184
rect 3762 2128 3790 2184
rect 3950 2128 3978 2184
rect 4414 2128 4442 2184
rect 4546 2128 4574 2184
rect 5010 2128 5038 2184
rect 5198 2128 5226 2184
rect 5662 2128 5690 2184
rect 5794 2128 5822 2184
rect 6258 2128 6286 2184
rect 6446 2128 6474 2184
rect 6910 2128 6938 2184
rect 7042 2128 7070 2184
rect 7506 2128 7534 2184
rect 7694 2128 7722 2184
rect 8158 2128 8186 2184
rect 8290 2128 8318 2184
rect 8754 2128 8782 2184
rect 8942 2128 8970 2184
rect 9406 2128 9434 2184
rect 9538 2128 9566 2184
rect 10002 2128 10030 2184
rect 10190 2128 10218 2184
rect 10654 2128 10682 2184
rect 10786 2128 10814 2184
rect 11250 2128 11278 2184
rect 11438 2128 11466 2184
rect 11902 2128 11930 2184
rect 12034 2128 12062 2184
rect 12498 2128 12526 2184
rect 12686 2128 12714 2184
rect 13150 2128 13178 2184
rect 13282 2128 13310 2184
rect 13746 2128 13774 2184
rect 13934 2128 13962 2184
rect 14398 2128 14426 2184
rect 14530 2128 14558 2184
rect 14994 2128 15022 2184
rect 15182 2128 15210 2184
rect 15646 2128 15674 2184
rect 15778 2128 15806 2184
rect 16242 2128 16270 2184
rect 16430 2128 16458 2184
rect 16894 2128 16922 2184
rect 17026 2128 17054 2184
rect 17490 2128 17518 2184
rect 17678 2128 17706 2184
rect 18142 2128 18170 2184
rect 18274 2128 18302 2184
rect 18738 2128 18766 2184
rect 18926 2128 18954 2184
rect 19390 2128 19418 2184
rect 19522 2128 19550 2184
rect 19986 2128 20014 2184
rect 20174 2128 20202 2184
rect 20638 2128 20666 2184
rect 20770 2128 20798 2184
rect 21234 2128 21262 2184
rect 21422 2128 21450 2184
rect 21886 2128 21914 2184
rect 22018 2128 22046 2184
rect 22482 2128 22510 2184
rect 22670 2128 22698 2184
rect 23134 2128 23162 2184
rect 23266 2128 23294 2184
rect 23730 2128 23758 2184
rect 23918 2128 23946 2184
rect 24382 2128 24410 2184
rect 24514 2128 24542 2184
rect 24978 2128 25006 2184
rect 25166 2128 25194 2184
rect 25630 2128 25658 2184
rect 25762 2128 25790 2184
rect 26226 2128 26254 2184
rect 26414 2128 26442 2184
rect 26878 2128 26906 2184
rect 27010 2128 27038 2184
rect 27474 2128 27502 2184
rect 27662 2128 27690 2184
rect 28126 2128 28154 2184
rect 28258 2128 28286 2184
rect 28722 2128 28750 2184
rect 28910 2128 28938 2184
rect 29374 2128 29402 2184
rect 29506 2128 29534 2184
rect 29970 2128 29998 2184
rect 30158 2128 30186 2184
rect 30622 2128 30650 2184
rect 30754 2128 30782 2184
rect 31218 2128 31246 2184
rect 31406 2128 31434 2184
rect 31870 2128 31898 2184
rect 32002 2128 32030 2184
rect 32466 2128 32494 2184
rect 32654 2128 32682 2184
rect 33118 2128 33146 2184
rect 33250 2128 33278 2184
rect 33714 2128 33742 2184
rect 33902 2128 33930 2184
rect 34366 2128 34394 2184
rect 34498 2128 34526 2184
rect 34962 2128 34990 2184
rect 35150 2128 35178 2184
rect 35614 2128 35642 2184
rect 35746 2128 35774 2184
rect 36210 2128 36238 2184
rect 36398 2128 36426 2184
rect 36862 2128 36890 2184
rect 36994 2128 37022 2184
rect 37458 2128 37486 2184
rect 37646 2128 37674 2184
rect 38110 2128 38138 2184
rect 38242 2128 38270 2184
rect 38706 2128 38734 2184
rect 38894 2128 38922 2184
rect 39358 2128 39386 2184
rect 39490 2128 39518 2184
rect 39954 2128 39982 2184
rect 40142 2128 40170 2184
rect 40606 2128 40634 2184
rect 40738 2128 40766 2184
rect 41202 2128 41230 2184
rect 41390 2128 41418 2184
rect 41854 2128 41882 2184
rect 41986 2128 42014 2184
rect 42450 2128 42478 2184
rect 42638 2128 42666 2184
rect 43102 2128 43130 2184
rect 43234 2128 43262 2184
rect 43698 2128 43726 2184
rect 43886 2128 43914 2184
rect 44350 2128 44378 2184
rect 44482 2128 44510 2184
rect 44946 2128 44974 2184
rect 45134 2128 45162 2184
rect 45598 2128 45626 2184
rect 45730 2128 45758 2184
rect 46194 2128 46222 2184
rect 46382 2128 46410 2184
rect 46846 2128 46874 2184
rect 46978 2128 47006 2184
rect 47442 2128 47470 2184
rect 47630 2128 47658 2184
rect 48094 2128 48122 2184
rect 48226 2128 48254 2184
rect 48690 2128 48718 2184
rect 48878 2128 48906 2184
rect 49342 2128 49370 2184
rect 49474 2128 49502 2184
rect 49938 2128 49966 2184
rect 50126 2128 50154 2184
rect 50590 2128 50618 2184
rect 50722 2128 50750 2184
rect 51186 2128 51214 2184
rect 51374 2128 51402 2184
rect 51838 2128 51866 2184
rect 51970 2128 51998 2184
rect 52434 2128 52462 2184
rect 52622 2128 52650 2184
rect 53086 2128 53114 2184
rect 53218 2128 53246 2184
rect 53682 2128 53710 2184
rect 53870 2128 53898 2184
rect 54334 2128 54362 2184
rect 54466 2128 54494 2184
rect 54930 2128 54958 2184
rect 55118 2128 55146 2184
rect 55582 2128 55610 2184
rect 55714 2128 55742 2184
rect 56178 2128 56206 2184
rect 56366 2128 56394 2184
rect 56830 2128 56858 2184
rect 56962 2128 56990 2184
rect 57426 2128 57454 2184
rect 57614 2128 57642 2184
rect 58078 2128 58106 2184
rect 58210 2128 58238 2184
rect 58674 2128 58702 2184
rect 58862 2128 58890 2184
rect 59326 2128 59354 2184
rect 59458 2128 59486 2184
rect 59922 2128 59950 2184
rect 60110 2128 60138 2184
rect 60574 2128 60602 2184
rect 60706 2128 60734 2184
rect 61170 2128 61198 2184
rect 61358 2128 61386 2184
rect 61822 2128 61850 2184
rect 61954 2128 61982 2184
rect 62418 2128 62446 2184
rect 62606 2128 62634 2184
rect 63070 2128 63098 2184
rect 63202 2128 63230 2184
rect 63666 2128 63694 2184
rect 63854 2128 63882 2184
rect 64318 2128 64346 2184
rect 64450 2128 64478 2184
rect 64914 2128 64942 2184
rect 65102 2128 65130 2184
rect 65566 2128 65594 2184
rect 65698 2128 65726 2184
rect 66162 2128 66190 2184
rect 66350 2128 66378 2184
rect 66814 2128 66842 2184
rect 66946 2128 66974 2184
rect 67410 2128 67438 2184
rect 67598 2128 67626 2184
rect 68062 2128 68090 2184
rect 68194 2128 68222 2184
rect 68658 2128 68686 2184
rect 68846 2128 68874 2184
rect 69310 2128 69338 2184
rect 69442 2128 69470 2184
rect 69906 2128 69934 2184
rect 70094 2128 70122 2184
rect 70558 2128 70586 2184
rect 70690 2128 70718 2184
rect 71154 2128 71182 2184
rect 71342 2128 71370 2184
rect 71806 2128 71834 2184
rect 71938 2128 71966 2184
rect 72402 2128 72430 2184
rect 72590 2128 72618 2184
rect 73054 2128 73082 2184
rect 73186 2128 73214 2184
rect 73650 2128 73678 2184
rect 73838 2128 73866 2184
rect 74302 2128 74330 2184
rect 74434 2128 74462 2184
rect 74898 2128 74926 2184
rect 75086 2128 75114 2184
rect 75550 2128 75578 2184
rect 75682 2128 75710 2184
rect 76146 2128 76174 2184
rect 76334 2128 76362 2184
rect 76798 2128 76826 2184
rect 76930 2128 76958 2184
rect 77394 2128 77422 2184
rect 77582 2128 77610 2184
rect 78046 2128 78074 2184
rect 78178 2128 78206 2184
rect 78642 2128 78670 2184
rect 78830 2128 78858 2184
rect 79294 2128 79322 2184
rect 79426 2128 79454 2184
rect 79890 2128 79918 2184
rect 80078 2128 80106 2184
rect 80542 2128 80570 2184
rect 80674 2128 80702 2184
rect 81138 2128 81166 2184
rect 1454 274 1482 868
rect 1654 376 1660 428
rect 1712 376 1718 428
rect 1436 222 1442 274
rect 1494 222 1500 274
rect 1918 150 1946 868
rect 2050 150 2078 868
rect 2278 500 2284 552
rect 2336 500 2342 552
rect 2514 274 2542 868
rect 2702 274 2730 868
rect 2902 624 2908 676
rect 2960 624 2966 676
rect 2496 222 2502 274
rect 2554 222 2560 274
rect 2684 222 2690 274
rect 2742 222 2748 274
rect 3166 150 3194 868
rect 3298 150 3326 868
rect 3526 748 3532 800
rect 3584 748 3590 800
rect 3762 274 3790 868
rect 3950 274 3978 868
rect 4150 376 4156 428
rect 4208 376 4214 428
rect 3744 222 3750 274
rect 3802 222 3808 274
rect 3932 222 3938 274
rect 3990 222 3996 274
rect 4414 150 4442 868
rect 4546 150 4574 868
rect 4774 500 4780 552
rect 4832 500 4838 552
rect 5010 274 5038 868
rect 5198 274 5226 868
rect 5398 624 5404 676
rect 5456 624 5462 676
rect 4992 222 4998 274
rect 5050 222 5056 274
rect 5180 222 5186 274
rect 5238 222 5244 274
rect 5662 150 5690 868
rect 5794 150 5822 868
rect 6022 748 6028 800
rect 6080 748 6086 800
rect 6258 274 6286 868
rect 6446 274 6474 868
rect 6646 376 6652 428
rect 6704 376 6710 428
rect 6240 222 6246 274
rect 6298 222 6304 274
rect 6428 222 6434 274
rect 6486 222 6492 274
rect 6910 150 6938 868
rect 7042 150 7070 868
rect 7270 500 7276 552
rect 7328 500 7334 552
rect 7506 274 7534 868
rect 7694 274 7722 868
rect 7894 624 7900 676
rect 7952 624 7958 676
rect 7488 222 7494 274
rect 7546 222 7552 274
rect 7676 222 7682 274
rect 7734 222 7740 274
rect 8158 150 8186 868
rect 8290 150 8318 868
rect 8518 748 8524 800
rect 8576 748 8582 800
rect 8754 274 8782 868
rect 8942 274 8970 868
rect 9142 376 9148 428
rect 9200 376 9206 428
rect 8736 222 8742 274
rect 8794 222 8800 274
rect 8924 222 8930 274
rect 8982 222 8988 274
rect 9406 150 9434 868
rect 9538 150 9566 868
rect 9766 500 9772 552
rect 9824 500 9830 552
rect 10002 274 10030 868
rect 10190 274 10218 868
rect 10390 624 10396 676
rect 10448 624 10454 676
rect 9984 222 9990 274
rect 10042 222 10048 274
rect 10172 222 10178 274
rect 10230 222 10236 274
rect 10654 150 10682 868
rect 10786 150 10814 868
rect 11014 748 11020 800
rect 11072 748 11078 800
rect 11250 274 11278 868
rect 11438 274 11466 868
rect 11638 376 11644 428
rect 11696 376 11702 428
rect 11232 222 11238 274
rect 11290 222 11296 274
rect 11420 222 11426 274
rect 11478 222 11484 274
rect 11902 150 11930 868
rect 12034 150 12062 868
rect 12262 500 12268 552
rect 12320 500 12326 552
rect 12498 274 12526 868
rect 12686 274 12714 868
rect 12886 624 12892 676
rect 12944 624 12950 676
rect 12480 222 12486 274
rect 12538 222 12544 274
rect 12668 222 12674 274
rect 12726 222 12732 274
rect 13150 150 13178 868
rect 13282 150 13310 868
rect 13510 748 13516 800
rect 13568 748 13574 800
rect 13746 274 13774 868
rect 13934 274 13962 868
rect 14134 376 14140 428
rect 14192 376 14198 428
rect 13728 222 13734 274
rect 13786 222 13792 274
rect 13916 222 13922 274
rect 13974 222 13980 274
rect 14398 150 14426 868
rect 14530 150 14558 868
rect 14758 500 14764 552
rect 14816 500 14822 552
rect 14994 274 15022 868
rect 15182 274 15210 868
rect 15382 624 15388 676
rect 15440 624 15446 676
rect 14976 222 14982 274
rect 15034 222 15040 274
rect 15164 222 15170 274
rect 15222 222 15228 274
rect 15646 150 15674 868
rect 15778 150 15806 868
rect 16006 748 16012 800
rect 16064 748 16070 800
rect 16242 274 16270 868
rect 16430 274 16458 868
rect 16630 376 16636 428
rect 16688 376 16694 428
rect 16224 222 16230 274
rect 16282 222 16288 274
rect 16412 222 16418 274
rect 16470 222 16476 274
rect 16894 150 16922 868
rect 17026 150 17054 868
rect 17254 500 17260 552
rect 17312 500 17318 552
rect 17490 274 17518 868
rect 17678 274 17706 868
rect 17878 624 17884 676
rect 17936 624 17942 676
rect 17472 222 17478 274
rect 17530 222 17536 274
rect 17660 222 17666 274
rect 17718 222 17724 274
rect 18142 150 18170 868
rect 18274 150 18302 868
rect 18502 748 18508 800
rect 18560 748 18566 800
rect 18738 274 18766 868
rect 18926 274 18954 868
rect 19126 376 19132 428
rect 19184 376 19190 428
rect 18720 222 18726 274
rect 18778 222 18784 274
rect 18908 222 18914 274
rect 18966 222 18972 274
rect 19390 150 19418 868
rect 19522 150 19550 868
rect 19750 500 19756 552
rect 19808 500 19814 552
rect 19986 274 20014 868
rect 20174 274 20202 868
rect 20374 624 20380 676
rect 20432 624 20438 676
rect 19968 222 19974 274
rect 20026 222 20032 274
rect 20156 222 20162 274
rect 20214 222 20220 274
rect 20638 150 20666 868
rect 20770 150 20798 868
rect 20998 748 21004 800
rect 21056 748 21062 800
rect 21234 274 21262 868
rect 21422 274 21450 868
rect 21622 376 21628 428
rect 21680 376 21686 428
rect 21216 222 21222 274
rect 21274 222 21280 274
rect 21404 222 21410 274
rect 21462 222 21468 274
rect 21886 150 21914 868
rect 22018 150 22046 868
rect 22246 500 22252 552
rect 22304 500 22310 552
rect 22482 274 22510 868
rect 22670 274 22698 868
rect 22870 624 22876 676
rect 22928 624 22934 676
rect 22464 222 22470 274
rect 22522 222 22528 274
rect 22652 222 22658 274
rect 22710 222 22716 274
rect 23134 150 23162 868
rect 23266 150 23294 868
rect 23494 748 23500 800
rect 23552 748 23558 800
rect 23730 274 23758 868
rect 23918 274 23946 868
rect 24118 376 24124 428
rect 24176 376 24182 428
rect 23712 222 23718 274
rect 23770 222 23776 274
rect 23900 222 23906 274
rect 23958 222 23964 274
rect 24382 150 24410 868
rect 24514 150 24542 868
rect 24742 500 24748 552
rect 24800 500 24806 552
rect 24978 274 25006 868
rect 25166 274 25194 868
rect 25366 624 25372 676
rect 25424 624 25430 676
rect 24960 222 24966 274
rect 25018 222 25024 274
rect 25148 222 25154 274
rect 25206 222 25212 274
rect 25630 150 25658 868
rect 25762 150 25790 868
rect 25990 748 25996 800
rect 26048 748 26054 800
rect 26226 274 26254 868
rect 26414 274 26442 868
rect 26614 376 26620 428
rect 26672 376 26678 428
rect 26208 222 26214 274
rect 26266 222 26272 274
rect 26396 222 26402 274
rect 26454 222 26460 274
rect 26878 150 26906 868
rect 27010 150 27038 868
rect 27238 500 27244 552
rect 27296 500 27302 552
rect 27474 274 27502 868
rect 27662 274 27690 868
rect 27862 624 27868 676
rect 27920 624 27926 676
rect 27456 222 27462 274
rect 27514 222 27520 274
rect 27644 222 27650 274
rect 27702 222 27708 274
rect 28126 150 28154 868
rect 28258 150 28286 868
rect 28486 748 28492 800
rect 28544 748 28550 800
rect 28722 274 28750 868
rect 28910 274 28938 868
rect 29110 376 29116 428
rect 29168 376 29174 428
rect 28704 222 28710 274
rect 28762 222 28768 274
rect 28892 222 28898 274
rect 28950 222 28956 274
rect 29374 150 29402 868
rect 29506 150 29534 868
rect 29734 500 29740 552
rect 29792 500 29798 552
rect 29970 274 29998 868
rect 30158 274 30186 868
rect 30358 624 30364 676
rect 30416 624 30422 676
rect 29952 222 29958 274
rect 30010 222 30016 274
rect 30140 222 30146 274
rect 30198 222 30204 274
rect 30622 150 30650 868
rect 30754 150 30782 868
rect 30982 748 30988 800
rect 31040 748 31046 800
rect 31218 274 31246 868
rect 31406 274 31434 868
rect 31606 376 31612 428
rect 31664 376 31670 428
rect 31200 222 31206 274
rect 31258 222 31264 274
rect 31388 222 31394 274
rect 31446 222 31452 274
rect 31870 150 31898 868
rect 32002 150 32030 868
rect 32230 500 32236 552
rect 32288 500 32294 552
rect 32466 274 32494 868
rect 32654 274 32682 868
rect 32854 624 32860 676
rect 32912 624 32918 676
rect 32448 222 32454 274
rect 32506 222 32512 274
rect 32636 222 32642 274
rect 32694 222 32700 274
rect 33118 150 33146 868
rect 33250 150 33278 868
rect 33478 748 33484 800
rect 33536 748 33542 800
rect 33714 274 33742 868
rect 33902 274 33930 868
rect 34102 376 34108 428
rect 34160 376 34166 428
rect 33696 222 33702 274
rect 33754 222 33760 274
rect 33884 222 33890 274
rect 33942 222 33948 274
rect 34366 150 34394 868
rect 34498 150 34526 868
rect 34726 500 34732 552
rect 34784 500 34790 552
rect 34962 274 34990 868
rect 35150 274 35178 868
rect 35350 624 35356 676
rect 35408 624 35414 676
rect 34944 222 34950 274
rect 35002 222 35008 274
rect 35132 222 35138 274
rect 35190 222 35196 274
rect 35614 150 35642 868
rect 35746 150 35774 868
rect 35974 748 35980 800
rect 36032 748 36038 800
rect 36210 274 36238 868
rect 36398 274 36426 868
rect 36598 376 36604 428
rect 36656 376 36662 428
rect 36192 222 36198 274
rect 36250 222 36256 274
rect 36380 222 36386 274
rect 36438 222 36444 274
rect 36862 150 36890 868
rect 36994 150 37022 868
rect 37222 500 37228 552
rect 37280 500 37286 552
rect 37458 274 37486 868
rect 37646 274 37674 868
rect 37846 624 37852 676
rect 37904 624 37910 676
rect 37440 222 37446 274
rect 37498 222 37504 274
rect 37628 222 37634 274
rect 37686 222 37692 274
rect 38110 150 38138 868
rect 38242 150 38270 868
rect 38470 748 38476 800
rect 38528 748 38534 800
rect 38706 274 38734 868
rect 38894 274 38922 868
rect 39094 376 39100 428
rect 39152 376 39158 428
rect 38688 222 38694 274
rect 38746 222 38752 274
rect 38876 222 38882 274
rect 38934 222 38940 274
rect 39358 150 39386 868
rect 39490 150 39518 868
rect 39718 500 39724 552
rect 39776 500 39782 552
rect 39954 274 39982 868
rect 40142 274 40170 868
rect 40342 624 40348 676
rect 40400 624 40406 676
rect 39936 222 39942 274
rect 39994 222 40000 274
rect 40124 222 40130 274
rect 40182 222 40188 274
rect 40606 150 40634 868
rect 40738 150 40766 868
rect 40966 748 40972 800
rect 41024 748 41030 800
rect 41202 274 41230 868
rect 41390 274 41418 868
rect 41590 376 41596 428
rect 41648 376 41654 428
rect 41184 222 41190 274
rect 41242 222 41248 274
rect 41372 222 41378 274
rect 41430 222 41436 274
rect 41854 150 41882 868
rect 41986 150 42014 868
rect 42214 500 42220 552
rect 42272 500 42278 552
rect 42450 274 42478 868
rect 42638 274 42666 868
rect 42838 624 42844 676
rect 42896 624 42902 676
rect 42432 222 42438 274
rect 42490 222 42496 274
rect 42620 222 42626 274
rect 42678 222 42684 274
rect 43102 150 43130 868
rect 43234 150 43262 868
rect 43462 748 43468 800
rect 43520 748 43526 800
rect 43698 274 43726 868
rect 43886 274 43914 868
rect 44086 376 44092 428
rect 44144 376 44150 428
rect 43680 222 43686 274
rect 43738 222 43744 274
rect 43868 222 43874 274
rect 43926 222 43932 274
rect 44350 150 44378 868
rect 44482 150 44510 868
rect 44710 500 44716 552
rect 44768 500 44774 552
rect 44946 274 44974 868
rect 45134 274 45162 868
rect 45334 624 45340 676
rect 45392 624 45398 676
rect 44928 222 44934 274
rect 44986 222 44992 274
rect 45116 222 45122 274
rect 45174 222 45180 274
rect 45598 150 45626 868
rect 45730 150 45758 868
rect 45958 748 45964 800
rect 46016 748 46022 800
rect 46194 274 46222 868
rect 46382 274 46410 868
rect 46582 376 46588 428
rect 46640 376 46646 428
rect 46176 222 46182 274
rect 46234 222 46240 274
rect 46364 222 46370 274
rect 46422 222 46428 274
rect 46846 150 46874 868
rect 46978 150 47006 868
rect 47206 500 47212 552
rect 47264 500 47270 552
rect 47442 274 47470 868
rect 47630 274 47658 868
rect 47830 624 47836 676
rect 47888 624 47894 676
rect 47424 222 47430 274
rect 47482 222 47488 274
rect 47612 222 47618 274
rect 47670 222 47676 274
rect 48094 150 48122 868
rect 48226 150 48254 868
rect 48454 748 48460 800
rect 48512 748 48518 800
rect 48690 274 48718 868
rect 48878 274 48906 868
rect 49078 376 49084 428
rect 49136 376 49142 428
rect 48672 222 48678 274
rect 48730 222 48736 274
rect 48860 222 48866 274
rect 48918 222 48924 274
rect 49342 150 49370 868
rect 49474 150 49502 868
rect 49702 500 49708 552
rect 49760 500 49766 552
rect 49938 274 49966 868
rect 50126 274 50154 868
rect 50326 624 50332 676
rect 50384 624 50390 676
rect 49920 222 49926 274
rect 49978 222 49984 274
rect 50108 222 50114 274
rect 50166 222 50172 274
rect 50590 150 50618 868
rect 50722 150 50750 868
rect 50950 748 50956 800
rect 51008 748 51014 800
rect 51186 274 51214 868
rect 51374 274 51402 868
rect 51574 376 51580 428
rect 51632 376 51638 428
rect 51168 222 51174 274
rect 51226 222 51232 274
rect 51356 222 51362 274
rect 51414 222 51420 274
rect 51838 150 51866 868
rect 51970 150 51998 868
rect 52198 500 52204 552
rect 52256 500 52262 552
rect 52434 274 52462 868
rect 52622 274 52650 868
rect 52822 624 52828 676
rect 52880 624 52886 676
rect 52416 222 52422 274
rect 52474 222 52480 274
rect 52604 222 52610 274
rect 52662 222 52668 274
rect 53086 150 53114 868
rect 53218 150 53246 868
rect 53446 748 53452 800
rect 53504 748 53510 800
rect 53682 274 53710 868
rect 53870 274 53898 868
rect 54070 376 54076 428
rect 54128 376 54134 428
rect 53664 222 53670 274
rect 53722 222 53728 274
rect 53852 222 53858 274
rect 53910 222 53916 274
rect 54334 150 54362 868
rect 54466 150 54494 868
rect 54694 500 54700 552
rect 54752 500 54758 552
rect 54930 274 54958 868
rect 55118 274 55146 868
rect 55318 624 55324 676
rect 55376 624 55382 676
rect 54912 222 54918 274
rect 54970 222 54976 274
rect 55100 222 55106 274
rect 55158 222 55164 274
rect 55582 150 55610 868
rect 55714 150 55742 868
rect 55942 748 55948 800
rect 56000 748 56006 800
rect 56178 274 56206 868
rect 56366 274 56394 868
rect 56566 376 56572 428
rect 56624 376 56630 428
rect 56160 222 56166 274
rect 56218 222 56224 274
rect 56348 222 56354 274
rect 56406 222 56412 274
rect 56830 150 56858 868
rect 56962 150 56990 868
rect 57190 500 57196 552
rect 57248 500 57254 552
rect 57426 274 57454 868
rect 57614 274 57642 868
rect 57814 624 57820 676
rect 57872 624 57878 676
rect 57408 222 57414 274
rect 57466 222 57472 274
rect 57596 222 57602 274
rect 57654 222 57660 274
rect 58078 150 58106 868
rect 58210 150 58238 868
rect 58438 748 58444 800
rect 58496 748 58502 800
rect 58674 274 58702 868
rect 58862 274 58890 868
rect 59062 376 59068 428
rect 59120 376 59126 428
rect 58656 222 58662 274
rect 58714 222 58720 274
rect 58844 222 58850 274
rect 58902 222 58908 274
rect 59326 150 59354 868
rect 59458 150 59486 868
rect 59686 500 59692 552
rect 59744 500 59750 552
rect 59922 274 59950 868
rect 60110 274 60138 868
rect 60310 624 60316 676
rect 60368 624 60374 676
rect 59904 222 59910 274
rect 59962 222 59968 274
rect 60092 222 60098 274
rect 60150 222 60156 274
rect 60574 150 60602 868
rect 60706 150 60734 868
rect 60934 748 60940 800
rect 60992 748 60998 800
rect 61170 274 61198 868
rect 61358 274 61386 868
rect 61558 376 61564 428
rect 61616 376 61622 428
rect 61152 222 61158 274
rect 61210 222 61216 274
rect 61340 222 61346 274
rect 61398 222 61404 274
rect 61822 150 61850 868
rect 61954 150 61982 868
rect 62182 500 62188 552
rect 62240 500 62246 552
rect 62418 274 62446 868
rect 62606 274 62634 868
rect 62806 624 62812 676
rect 62864 624 62870 676
rect 62400 222 62406 274
rect 62458 222 62464 274
rect 62588 222 62594 274
rect 62646 222 62652 274
rect 63070 150 63098 868
rect 63202 150 63230 868
rect 63430 748 63436 800
rect 63488 748 63494 800
rect 63666 274 63694 868
rect 63854 274 63882 868
rect 64054 376 64060 428
rect 64112 376 64118 428
rect 63648 222 63654 274
rect 63706 222 63712 274
rect 63836 222 63842 274
rect 63894 222 63900 274
rect 64318 150 64346 868
rect 64450 150 64478 868
rect 64678 500 64684 552
rect 64736 500 64742 552
rect 64914 274 64942 868
rect 65102 274 65130 868
rect 65302 624 65308 676
rect 65360 624 65366 676
rect 64896 222 64902 274
rect 64954 222 64960 274
rect 65084 222 65090 274
rect 65142 222 65148 274
rect 65566 150 65594 868
rect 65698 150 65726 868
rect 65926 748 65932 800
rect 65984 748 65990 800
rect 66162 274 66190 868
rect 66350 274 66378 868
rect 66550 376 66556 428
rect 66608 376 66614 428
rect 66144 222 66150 274
rect 66202 222 66208 274
rect 66332 222 66338 274
rect 66390 222 66396 274
rect 66814 150 66842 868
rect 66946 150 66974 868
rect 67174 500 67180 552
rect 67232 500 67238 552
rect 67410 274 67438 868
rect 67598 274 67626 868
rect 67798 624 67804 676
rect 67856 624 67862 676
rect 67392 222 67398 274
rect 67450 222 67456 274
rect 67580 222 67586 274
rect 67638 222 67644 274
rect 68062 150 68090 868
rect 68194 150 68222 868
rect 68422 748 68428 800
rect 68480 748 68486 800
rect 68658 274 68686 868
rect 68846 274 68874 868
rect 69046 376 69052 428
rect 69104 376 69110 428
rect 68640 222 68646 274
rect 68698 222 68704 274
rect 68828 222 68834 274
rect 68886 222 68892 274
rect 69310 150 69338 868
rect 69442 150 69470 868
rect 69670 500 69676 552
rect 69728 500 69734 552
rect 69906 274 69934 868
rect 70094 274 70122 868
rect 70294 624 70300 676
rect 70352 624 70358 676
rect 69888 222 69894 274
rect 69946 222 69952 274
rect 70076 222 70082 274
rect 70134 222 70140 274
rect 70558 150 70586 868
rect 70690 150 70718 868
rect 70918 748 70924 800
rect 70976 748 70982 800
rect 71154 274 71182 868
rect 71342 274 71370 868
rect 71542 376 71548 428
rect 71600 376 71606 428
rect 71136 222 71142 274
rect 71194 222 71200 274
rect 71324 222 71330 274
rect 71382 222 71388 274
rect 71806 150 71834 868
rect 71938 150 71966 868
rect 72166 500 72172 552
rect 72224 500 72230 552
rect 72402 274 72430 868
rect 72590 274 72618 868
rect 72790 624 72796 676
rect 72848 624 72854 676
rect 72384 222 72390 274
rect 72442 222 72448 274
rect 72572 222 72578 274
rect 72630 222 72636 274
rect 73054 150 73082 868
rect 73186 150 73214 868
rect 73414 748 73420 800
rect 73472 748 73478 800
rect 73650 274 73678 868
rect 73838 274 73866 868
rect 74038 376 74044 428
rect 74096 376 74102 428
rect 73632 222 73638 274
rect 73690 222 73696 274
rect 73820 222 73826 274
rect 73878 222 73884 274
rect 74302 150 74330 868
rect 74434 150 74462 868
rect 74662 500 74668 552
rect 74720 500 74726 552
rect 74898 274 74926 868
rect 75086 274 75114 868
rect 75286 624 75292 676
rect 75344 624 75350 676
rect 74880 222 74886 274
rect 74938 222 74944 274
rect 75068 222 75074 274
rect 75126 222 75132 274
rect 75550 150 75578 868
rect 75682 150 75710 868
rect 75910 748 75916 800
rect 75968 748 75974 800
rect 76146 274 76174 868
rect 76334 274 76362 868
rect 76534 376 76540 428
rect 76592 376 76598 428
rect 76128 222 76134 274
rect 76186 222 76192 274
rect 76316 222 76322 274
rect 76374 222 76380 274
rect 76798 150 76826 868
rect 76930 150 76958 868
rect 77158 500 77164 552
rect 77216 500 77222 552
rect 77394 274 77422 868
rect 77582 274 77610 868
rect 77782 624 77788 676
rect 77840 624 77846 676
rect 77376 222 77382 274
rect 77434 222 77440 274
rect 77564 222 77570 274
rect 77622 222 77628 274
rect 78046 150 78074 868
rect 78178 150 78206 868
rect 78406 748 78412 800
rect 78464 748 78470 800
rect 78642 274 78670 868
rect 78830 274 78858 868
rect 79030 376 79036 428
rect 79088 376 79094 428
rect 78624 222 78630 274
rect 78682 222 78688 274
rect 78812 222 78818 274
rect 78870 222 78876 274
rect 79294 150 79322 868
rect 79426 150 79454 868
rect 79654 500 79660 552
rect 79712 500 79718 552
rect 79890 274 79918 868
rect 80078 274 80106 868
rect 80278 624 80284 676
rect 80336 624 80342 676
rect 79872 222 79878 274
rect 79930 222 79936 274
rect 80060 222 80066 274
rect 80118 222 80124 274
rect 80542 150 80570 868
rect 80674 150 80702 868
rect 80902 748 80908 800
rect 80960 748 80966 800
rect 81138 274 81166 868
rect 81120 222 81126 274
rect 81178 222 81184 274
rect 1900 98 1906 150
rect 1958 98 1964 150
rect 2032 98 2038 150
rect 2090 98 2096 150
rect 3148 98 3154 150
rect 3206 98 3212 150
rect 3280 98 3286 150
rect 3338 98 3344 150
rect 4396 98 4402 150
rect 4454 98 4460 150
rect 4528 98 4534 150
rect 4586 98 4592 150
rect 5644 98 5650 150
rect 5702 98 5708 150
rect 5776 98 5782 150
rect 5834 98 5840 150
rect 6892 98 6898 150
rect 6950 98 6956 150
rect 7024 98 7030 150
rect 7082 98 7088 150
rect 8140 98 8146 150
rect 8198 98 8204 150
rect 8272 98 8278 150
rect 8330 98 8336 150
rect 9388 98 9394 150
rect 9446 98 9452 150
rect 9520 98 9526 150
rect 9578 98 9584 150
rect 10636 98 10642 150
rect 10694 98 10700 150
rect 10768 98 10774 150
rect 10826 98 10832 150
rect 11884 98 11890 150
rect 11942 98 11948 150
rect 12016 98 12022 150
rect 12074 98 12080 150
rect 13132 98 13138 150
rect 13190 98 13196 150
rect 13264 98 13270 150
rect 13322 98 13328 150
rect 14380 98 14386 150
rect 14438 98 14444 150
rect 14512 98 14518 150
rect 14570 98 14576 150
rect 15628 98 15634 150
rect 15686 98 15692 150
rect 15760 98 15766 150
rect 15818 98 15824 150
rect 16876 98 16882 150
rect 16934 98 16940 150
rect 17008 98 17014 150
rect 17066 98 17072 150
rect 18124 98 18130 150
rect 18182 98 18188 150
rect 18256 98 18262 150
rect 18314 98 18320 150
rect 19372 98 19378 150
rect 19430 98 19436 150
rect 19504 98 19510 150
rect 19562 98 19568 150
rect 20620 98 20626 150
rect 20678 98 20684 150
rect 20752 98 20758 150
rect 20810 98 20816 150
rect 21868 98 21874 150
rect 21926 98 21932 150
rect 22000 98 22006 150
rect 22058 98 22064 150
rect 23116 98 23122 150
rect 23174 98 23180 150
rect 23248 98 23254 150
rect 23306 98 23312 150
rect 24364 98 24370 150
rect 24422 98 24428 150
rect 24496 98 24502 150
rect 24554 98 24560 150
rect 25612 98 25618 150
rect 25670 98 25676 150
rect 25744 98 25750 150
rect 25802 98 25808 150
rect 26860 98 26866 150
rect 26918 98 26924 150
rect 26992 98 26998 150
rect 27050 98 27056 150
rect 28108 98 28114 150
rect 28166 98 28172 150
rect 28240 98 28246 150
rect 28298 98 28304 150
rect 29356 98 29362 150
rect 29414 98 29420 150
rect 29488 98 29494 150
rect 29546 98 29552 150
rect 30604 98 30610 150
rect 30662 98 30668 150
rect 30736 98 30742 150
rect 30794 98 30800 150
rect 31852 98 31858 150
rect 31910 98 31916 150
rect 31984 98 31990 150
rect 32042 98 32048 150
rect 33100 98 33106 150
rect 33158 98 33164 150
rect 33232 98 33238 150
rect 33290 98 33296 150
rect 34348 98 34354 150
rect 34406 98 34412 150
rect 34480 98 34486 150
rect 34538 98 34544 150
rect 35596 98 35602 150
rect 35654 98 35660 150
rect 35728 98 35734 150
rect 35786 98 35792 150
rect 36844 98 36850 150
rect 36902 98 36908 150
rect 36976 98 36982 150
rect 37034 98 37040 150
rect 38092 98 38098 150
rect 38150 98 38156 150
rect 38224 98 38230 150
rect 38282 98 38288 150
rect 39340 98 39346 150
rect 39398 98 39404 150
rect 39472 98 39478 150
rect 39530 98 39536 150
rect 40588 98 40594 150
rect 40646 98 40652 150
rect 40720 98 40726 150
rect 40778 98 40784 150
rect 41836 98 41842 150
rect 41894 98 41900 150
rect 41968 98 41974 150
rect 42026 98 42032 150
rect 43084 98 43090 150
rect 43142 98 43148 150
rect 43216 98 43222 150
rect 43274 98 43280 150
rect 44332 98 44338 150
rect 44390 98 44396 150
rect 44464 98 44470 150
rect 44522 98 44528 150
rect 45580 98 45586 150
rect 45638 98 45644 150
rect 45712 98 45718 150
rect 45770 98 45776 150
rect 46828 98 46834 150
rect 46886 98 46892 150
rect 46960 98 46966 150
rect 47018 98 47024 150
rect 48076 98 48082 150
rect 48134 98 48140 150
rect 48208 98 48214 150
rect 48266 98 48272 150
rect 49324 98 49330 150
rect 49382 98 49388 150
rect 49456 98 49462 150
rect 49514 98 49520 150
rect 50572 98 50578 150
rect 50630 98 50636 150
rect 50704 98 50710 150
rect 50762 98 50768 150
rect 51820 98 51826 150
rect 51878 98 51884 150
rect 51952 98 51958 150
rect 52010 98 52016 150
rect 53068 98 53074 150
rect 53126 98 53132 150
rect 53200 98 53206 150
rect 53258 98 53264 150
rect 54316 98 54322 150
rect 54374 98 54380 150
rect 54448 98 54454 150
rect 54506 98 54512 150
rect 55564 98 55570 150
rect 55622 98 55628 150
rect 55696 98 55702 150
rect 55754 98 55760 150
rect 56812 98 56818 150
rect 56870 98 56876 150
rect 56944 98 56950 150
rect 57002 98 57008 150
rect 58060 98 58066 150
rect 58118 98 58124 150
rect 58192 98 58198 150
rect 58250 98 58256 150
rect 59308 98 59314 150
rect 59366 98 59372 150
rect 59440 98 59446 150
rect 59498 98 59504 150
rect 60556 98 60562 150
rect 60614 98 60620 150
rect 60688 98 60694 150
rect 60746 98 60752 150
rect 61804 98 61810 150
rect 61862 98 61868 150
rect 61936 98 61942 150
rect 61994 98 62000 150
rect 63052 98 63058 150
rect 63110 98 63116 150
rect 63184 98 63190 150
rect 63242 98 63248 150
rect 64300 98 64306 150
rect 64358 98 64364 150
rect 64432 98 64438 150
rect 64490 98 64496 150
rect 65548 98 65554 150
rect 65606 98 65612 150
rect 65680 98 65686 150
rect 65738 98 65744 150
rect 66796 98 66802 150
rect 66854 98 66860 150
rect 66928 98 66934 150
rect 66986 98 66992 150
rect 68044 98 68050 150
rect 68102 98 68108 150
rect 68176 98 68182 150
rect 68234 98 68240 150
rect 69292 98 69298 150
rect 69350 98 69356 150
rect 69424 98 69430 150
rect 69482 98 69488 150
rect 70540 98 70546 150
rect 70598 98 70604 150
rect 70672 98 70678 150
rect 70730 98 70736 150
rect 71788 98 71794 150
rect 71846 98 71852 150
rect 71920 98 71926 150
rect 71978 98 71984 150
rect 73036 98 73042 150
rect 73094 98 73100 150
rect 73168 98 73174 150
rect 73226 98 73232 150
rect 74284 98 74290 150
rect 74342 98 74348 150
rect 74416 98 74422 150
rect 74474 98 74480 150
rect 75532 98 75538 150
rect 75590 98 75596 150
rect 75664 98 75670 150
rect 75722 98 75728 150
rect 76780 98 76786 150
rect 76838 98 76844 150
rect 76912 98 76918 150
rect 76970 98 76976 150
rect 78028 98 78034 150
rect 78086 98 78092 150
rect 78160 98 78166 150
rect 78218 98 78224 150
rect 79276 98 79282 150
rect 79334 98 79340 150
rect 79408 98 79414 150
rect 79466 98 79472 150
rect 80524 98 80530 150
rect 80582 98 80588 150
rect 80656 98 80662 150
rect 80714 98 80720 150
<< via1 >>
rect 1660 419 1712 428
rect 1660 385 1669 419
rect 1669 385 1703 419
rect 1703 385 1712 419
rect 1660 376 1712 385
rect 1442 222 1494 274
rect 2284 543 2336 552
rect 2284 509 2293 543
rect 2293 509 2327 543
rect 2327 509 2336 543
rect 2284 500 2336 509
rect 2908 667 2960 676
rect 2908 633 2917 667
rect 2917 633 2951 667
rect 2951 633 2960 667
rect 2908 624 2960 633
rect 2502 222 2554 274
rect 2690 222 2742 274
rect 3532 791 3584 800
rect 3532 757 3541 791
rect 3541 757 3575 791
rect 3575 757 3584 791
rect 3532 748 3584 757
rect 4156 419 4208 428
rect 4156 385 4165 419
rect 4165 385 4199 419
rect 4199 385 4208 419
rect 4156 376 4208 385
rect 3750 222 3802 274
rect 3938 222 3990 274
rect 4780 543 4832 552
rect 4780 509 4789 543
rect 4789 509 4823 543
rect 4823 509 4832 543
rect 4780 500 4832 509
rect 5404 667 5456 676
rect 5404 633 5413 667
rect 5413 633 5447 667
rect 5447 633 5456 667
rect 5404 624 5456 633
rect 4998 222 5050 274
rect 5186 222 5238 274
rect 6028 791 6080 800
rect 6028 757 6037 791
rect 6037 757 6071 791
rect 6071 757 6080 791
rect 6028 748 6080 757
rect 6652 419 6704 428
rect 6652 385 6661 419
rect 6661 385 6695 419
rect 6695 385 6704 419
rect 6652 376 6704 385
rect 6246 222 6298 274
rect 6434 222 6486 274
rect 7276 543 7328 552
rect 7276 509 7285 543
rect 7285 509 7319 543
rect 7319 509 7328 543
rect 7276 500 7328 509
rect 7900 667 7952 676
rect 7900 633 7909 667
rect 7909 633 7943 667
rect 7943 633 7952 667
rect 7900 624 7952 633
rect 7494 222 7546 274
rect 7682 222 7734 274
rect 8524 791 8576 800
rect 8524 757 8533 791
rect 8533 757 8567 791
rect 8567 757 8576 791
rect 8524 748 8576 757
rect 9148 419 9200 428
rect 9148 385 9157 419
rect 9157 385 9191 419
rect 9191 385 9200 419
rect 9148 376 9200 385
rect 8742 222 8794 274
rect 8930 222 8982 274
rect 9772 543 9824 552
rect 9772 509 9781 543
rect 9781 509 9815 543
rect 9815 509 9824 543
rect 9772 500 9824 509
rect 10396 667 10448 676
rect 10396 633 10405 667
rect 10405 633 10439 667
rect 10439 633 10448 667
rect 10396 624 10448 633
rect 9990 222 10042 274
rect 10178 222 10230 274
rect 11020 791 11072 800
rect 11020 757 11029 791
rect 11029 757 11063 791
rect 11063 757 11072 791
rect 11020 748 11072 757
rect 11644 419 11696 428
rect 11644 385 11653 419
rect 11653 385 11687 419
rect 11687 385 11696 419
rect 11644 376 11696 385
rect 11238 222 11290 274
rect 11426 222 11478 274
rect 12268 543 12320 552
rect 12268 509 12277 543
rect 12277 509 12311 543
rect 12311 509 12320 543
rect 12268 500 12320 509
rect 12892 667 12944 676
rect 12892 633 12901 667
rect 12901 633 12935 667
rect 12935 633 12944 667
rect 12892 624 12944 633
rect 12486 222 12538 274
rect 12674 222 12726 274
rect 13516 791 13568 800
rect 13516 757 13525 791
rect 13525 757 13559 791
rect 13559 757 13568 791
rect 13516 748 13568 757
rect 14140 419 14192 428
rect 14140 385 14149 419
rect 14149 385 14183 419
rect 14183 385 14192 419
rect 14140 376 14192 385
rect 13734 222 13786 274
rect 13922 222 13974 274
rect 14764 543 14816 552
rect 14764 509 14773 543
rect 14773 509 14807 543
rect 14807 509 14816 543
rect 14764 500 14816 509
rect 15388 667 15440 676
rect 15388 633 15397 667
rect 15397 633 15431 667
rect 15431 633 15440 667
rect 15388 624 15440 633
rect 14982 222 15034 274
rect 15170 222 15222 274
rect 16012 791 16064 800
rect 16012 757 16021 791
rect 16021 757 16055 791
rect 16055 757 16064 791
rect 16012 748 16064 757
rect 16636 419 16688 428
rect 16636 385 16645 419
rect 16645 385 16679 419
rect 16679 385 16688 419
rect 16636 376 16688 385
rect 16230 222 16282 274
rect 16418 222 16470 274
rect 17260 543 17312 552
rect 17260 509 17269 543
rect 17269 509 17303 543
rect 17303 509 17312 543
rect 17260 500 17312 509
rect 17884 667 17936 676
rect 17884 633 17893 667
rect 17893 633 17927 667
rect 17927 633 17936 667
rect 17884 624 17936 633
rect 17478 222 17530 274
rect 17666 222 17718 274
rect 18508 791 18560 800
rect 18508 757 18517 791
rect 18517 757 18551 791
rect 18551 757 18560 791
rect 18508 748 18560 757
rect 19132 419 19184 428
rect 19132 385 19141 419
rect 19141 385 19175 419
rect 19175 385 19184 419
rect 19132 376 19184 385
rect 18726 222 18778 274
rect 18914 222 18966 274
rect 19756 543 19808 552
rect 19756 509 19765 543
rect 19765 509 19799 543
rect 19799 509 19808 543
rect 19756 500 19808 509
rect 20380 667 20432 676
rect 20380 633 20389 667
rect 20389 633 20423 667
rect 20423 633 20432 667
rect 20380 624 20432 633
rect 19974 222 20026 274
rect 20162 222 20214 274
rect 21004 791 21056 800
rect 21004 757 21013 791
rect 21013 757 21047 791
rect 21047 757 21056 791
rect 21004 748 21056 757
rect 21628 419 21680 428
rect 21628 385 21637 419
rect 21637 385 21671 419
rect 21671 385 21680 419
rect 21628 376 21680 385
rect 21222 222 21274 274
rect 21410 222 21462 274
rect 22252 543 22304 552
rect 22252 509 22261 543
rect 22261 509 22295 543
rect 22295 509 22304 543
rect 22252 500 22304 509
rect 22876 667 22928 676
rect 22876 633 22885 667
rect 22885 633 22919 667
rect 22919 633 22928 667
rect 22876 624 22928 633
rect 22470 222 22522 274
rect 22658 222 22710 274
rect 23500 791 23552 800
rect 23500 757 23509 791
rect 23509 757 23543 791
rect 23543 757 23552 791
rect 23500 748 23552 757
rect 24124 419 24176 428
rect 24124 385 24133 419
rect 24133 385 24167 419
rect 24167 385 24176 419
rect 24124 376 24176 385
rect 23718 222 23770 274
rect 23906 222 23958 274
rect 24748 543 24800 552
rect 24748 509 24757 543
rect 24757 509 24791 543
rect 24791 509 24800 543
rect 24748 500 24800 509
rect 25372 667 25424 676
rect 25372 633 25381 667
rect 25381 633 25415 667
rect 25415 633 25424 667
rect 25372 624 25424 633
rect 24966 222 25018 274
rect 25154 222 25206 274
rect 25996 791 26048 800
rect 25996 757 26005 791
rect 26005 757 26039 791
rect 26039 757 26048 791
rect 25996 748 26048 757
rect 26620 419 26672 428
rect 26620 385 26629 419
rect 26629 385 26663 419
rect 26663 385 26672 419
rect 26620 376 26672 385
rect 26214 222 26266 274
rect 26402 222 26454 274
rect 27244 543 27296 552
rect 27244 509 27253 543
rect 27253 509 27287 543
rect 27287 509 27296 543
rect 27244 500 27296 509
rect 27868 667 27920 676
rect 27868 633 27877 667
rect 27877 633 27911 667
rect 27911 633 27920 667
rect 27868 624 27920 633
rect 27462 222 27514 274
rect 27650 222 27702 274
rect 28492 791 28544 800
rect 28492 757 28501 791
rect 28501 757 28535 791
rect 28535 757 28544 791
rect 28492 748 28544 757
rect 29116 419 29168 428
rect 29116 385 29125 419
rect 29125 385 29159 419
rect 29159 385 29168 419
rect 29116 376 29168 385
rect 28710 222 28762 274
rect 28898 222 28950 274
rect 29740 543 29792 552
rect 29740 509 29749 543
rect 29749 509 29783 543
rect 29783 509 29792 543
rect 29740 500 29792 509
rect 30364 667 30416 676
rect 30364 633 30373 667
rect 30373 633 30407 667
rect 30407 633 30416 667
rect 30364 624 30416 633
rect 29958 222 30010 274
rect 30146 222 30198 274
rect 30988 791 31040 800
rect 30988 757 30997 791
rect 30997 757 31031 791
rect 31031 757 31040 791
rect 30988 748 31040 757
rect 31612 419 31664 428
rect 31612 385 31621 419
rect 31621 385 31655 419
rect 31655 385 31664 419
rect 31612 376 31664 385
rect 31206 222 31258 274
rect 31394 222 31446 274
rect 32236 543 32288 552
rect 32236 509 32245 543
rect 32245 509 32279 543
rect 32279 509 32288 543
rect 32236 500 32288 509
rect 32860 667 32912 676
rect 32860 633 32869 667
rect 32869 633 32903 667
rect 32903 633 32912 667
rect 32860 624 32912 633
rect 32454 222 32506 274
rect 32642 222 32694 274
rect 33484 791 33536 800
rect 33484 757 33493 791
rect 33493 757 33527 791
rect 33527 757 33536 791
rect 33484 748 33536 757
rect 34108 419 34160 428
rect 34108 385 34117 419
rect 34117 385 34151 419
rect 34151 385 34160 419
rect 34108 376 34160 385
rect 33702 222 33754 274
rect 33890 222 33942 274
rect 34732 543 34784 552
rect 34732 509 34741 543
rect 34741 509 34775 543
rect 34775 509 34784 543
rect 34732 500 34784 509
rect 35356 667 35408 676
rect 35356 633 35365 667
rect 35365 633 35399 667
rect 35399 633 35408 667
rect 35356 624 35408 633
rect 34950 222 35002 274
rect 35138 222 35190 274
rect 35980 791 36032 800
rect 35980 757 35989 791
rect 35989 757 36023 791
rect 36023 757 36032 791
rect 35980 748 36032 757
rect 36604 419 36656 428
rect 36604 385 36613 419
rect 36613 385 36647 419
rect 36647 385 36656 419
rect 36604 376 36656 385
rect 36198 222 36250 274
rect 36386 222 36438 274
rect 37228 543 37280 552
rect 37228 509 37237 543
rect 37237 509 37271 543
rect 37271 509 37280 543
rect 37228 500 37280 509
rect 37852 667 37904 676
rect 37852 633 37861 667
rect 37861 633 37895 667
rect 37895 633 37904 667
rect 37852 624 37904 633
rect 37446 222 37498 274
rect 37634 222 37686 274
rect 38476 791 38528 800
rect 38476 757 38485 791
rect 38485 757 38519 791
rect 38519 757 38528 791
rect 38476 748 38528 757
rect 39100 419 39152 428
rect 39100 385 39109 419
rect 39109 385 39143 419
rect 39143 385 39152 419
rect 39100 376 39152 385
rect 38694 222 38746 274
rect 38882 222 38934 274
rect 39724 543 39776 552
rect 39724 509 39733 543
rect 39733 509 39767 543
rect 39767 509 39776 543
rect 39724 500 39776 509
rect 40348 667 40400 676
rect 40348 633 40357 667
rect 40357 633 40391 667
rect 40391 633 40400 667
rect 40348 624 40400 633
rect 39942 222 39994 274
rect 40130 222 40182 274
rect 40972 791 41024 800
rect 40972 757 40981 791
rect 40981 757 41015 791
rect 41015 757 41024 791
rect 40972 748 41024 757
rect 41596 419 41648 428
rect 41596 385 41605 419
rect 41605 385 41639 419
rect 41639 385 41648 419
rect 41596 376 41648 385
rect 41190 222 41242 274
rect 41378 222 41430 274
rect 42220 543 42272 552
rect 42220 509 42229 543
rect 42229 509 42263 543
rect 42263 509 42272 543
rect 42220 500 42272 509
rect 42844 667 42896 676
rect 42844 633 42853 667
rect 42853 633 42887 667
rect 42887 633 42896 667
rect 42844 624 42896 633
rect 42438 222 42490 274
rect 42626 222 42678 274
rect 43468 791 43520 800
rect 43468 757 43477 791
rect 43477 757 43511 791
rect 43511 757 43520 791
rect 43468 748 43520 757
rect 44092 419 44144 428
rect 44092 385 44101 419
rect 44101 385 44135 419
rect 44135 385 44144 419
rect 44092 376 44144 385
rect 43686 222 43738 274
rect 43874 222 43926 274
rect 44716 543 44768 552
rect 44716 509 44725 543
rect 44725 509 44759 543
rect 44759 509 44768 543
rect 44716 500 44768 509
rect 45340 667 45392 676
rect 45340 633 45349 667
rect 45349 633 45383 667
rect 45383 633 45392 667
rect 45340 624 45392 633
rect 44934 222 44986 274
rect 45122 222 45174 274
rect 45964 791 46016 800
rect 45964 757 45973 791
rect 45973 757 46007 791
rect 46007 757 46016 791
rect 45964 748 46016 757
rect 46588 419 46640 428
rect 46588 385 46597 419
rect 46597 385 46631 419
rect 46631 385 46640 419
rect 46588 376 46640 385
rect 46182 222 46234 274
rect 46370 222 46422 274
rect 47212 543 47264 552
rect 47212 509 47221 543
rect 47221 509 47255 543
rect 47255 509 47264 543
rect 47212 500 47264 509
rect 47836 667 47888 676
rect 47836 633 47845 667
rect 47845 633 47879 667
rect 47879 633 47888 667
rect 47836 624 47888 633
rect 47430 222 47482 274
rect 47618 222 47670 274
rect 48460 791 48512 800
rect 48460 757 48469 791
rect 48469 757 48503 791
rect 48503 757 48512 791
rect 48460 748 48512 757
rect 49084 419 49136 428
rect 49084 385 49093 419
rect 49093 385 49127 419
rect 49127 385 49136 419
rect 49084 376 49136 385
rect 48678 222 48730 274
rect 48866 222 48918 274
rect 49708 543 49760 552
rect 49708 509 49717 543
rect 49717 509 49751 543
rect 49751 509 49760 543
rect 49708 500 49760 509
rect 50332 667 50384 676
rect 50332 633 50341 667
rect 50341 633 50375 667
rect 50375 633 50384 667
rect 50332 624 50384 633
rect 49926 222 49978 274
rect 50114 222 50166 274
rect 50956 791 51008 800
rect 50956 757 50965 791
rect 50965 757 50999 791
rect 50999 757 51008 791
rect 50956 748 51008 757
rect 51580 419 51632 428
rect 51580 385 51589 419
rect 51589 385 51623 419
rect 51623 385 51632 419
rect 51580 376 51632 385
rect 51174 222 51226 274
rect 51362 222 51414 274
rect 52204 543 52256 552
rect 52204 509 52213 543
rect 52213 509 52247 543
rect 52247 509 52256 543
rect 52204 500 52256 509
rect 52828 667 52880 676
rect 52828 633 52837 667
rect 52837 633 52871 667
rect 52871 633 52880 667
rect 52828 624 52880 633
rect 52422 222 52474 274
rect 52610 222 52662 274
rect 53452 791 53504 800
rect 53452 757 53461 791
rect 53461 757 53495 791
rect 53495 757 53504 791
rect 53452 748 53504 757
rect 54076 419 54128 428
rect 54076 385 54085 419
rect 54085 385 54119 419
rect 54119 385 54128 419
rect 54076 376 54128 385
rect 53670 222 53722 274
rect 53858 222 53910 274
rect 54700 543 54752 552
rect 54700 509 54709 543
rect 54709 509 54743 543
rect 54743 509 54752 543
rect 54700 500 54752 509
rect 55324 667 55376 676
rect 55324 633 55333 667
rect 55333 633 55367 667
rect 55367 633 55376 667
rect 55324 624 55376 633
rect 54918 222 54970 274
rect 55106 222 55158 274
rect 55948 791 56000 800
rect 55948 757 55957 791
rect 55957 757 55991 791
rect 55991 757 56000 791
rect 55948 748 56000 757
rect 56572 419 56624 428
rect 56572 385 56581 419
rect 56581 385 56615 419
rect 56615 385 56624 419
rect 56572 376 56624 385
rect 56166 222 56218 274
rect 56354 222 56406 274
rect 57196 543 57248 552
rect 57196 509 57205 543
rect 57205 509 57239 543
rect 57239 509 57248 543
rect 57196 500 57248 509
rect 57820 667 57872 676
rect 57820 633 57829 667
rect 57829 633 57863 667
rect 57863 633 57872 667
rect 57820 624 57872 633
rect 57414 222 57466 274
rect 57602 222 57654 274
rect 58444 791 58496 800
rect 58444 757 58453 791
rect 58453 757 58487 791
rect 58487 757 58496 791
rect 58444 748 58496 757
rect 59068 419 59120 428
rect 59068 385 59077 419
rect 59077 385 59111 419
rect 59111 385 59120 419
rect 59068 376 59120 385
rect 58662 222 58714 274
rect 58850 222 58902 274
rect 59692 543 59744 552
rect 59692 509 59701 543
rect 59701 509 59735 543
rect 59735 509 59744 543
rect 59692 500 59744 509
rect 60316 667 60368 676
rect 60316 633 60325 667
rect 60325 633 60359 667
rect 60359 633 60368 667
rect 60316 624 60368 633
rect 59910 222 59962 274
rect 60098 222 60150 274
rect 60940 791 60992 800
rect 60940 757 60949 791
rect 60949 757 60983 791
rect 60983 757 60992 791
rect 60940 748 60992 757
rect 61564 419 61616 428
rect 61564 385 61573 419
rect 61573 385 61607 419
rect 61607 385 61616 419
rect 61564 376 61616 385
rect 61158 222 61210 274
rect 61346 222 61398 274
rect 62188 543 62240 552
rect 62188 509 62197 543
rect 62197 509 62231 543
rect 62231 509 62240 543
rect 62188 500 62240 509
rect 62812 667 62864 676
rect 62812 633 62821 667
rect 62821 633 62855 667
rect 62855 633 62864 667
rect 62812 624 62864 633
rect 62406 222 62458 274
rect 62594 222 62646 274
rect 63436 791 63488 800
rect 63436 757 63445 791
rect 63445 757 63479 791
rect 63479 757 63488 791
rect 63436 748 63488 757
rect 64060 419 64112 428
rect 64060 385 64069 419
rect 64069 385 64103 419
rect 64103 385 64112 419
rect 64060 376 64112 385
rect 63654 222 63706 274
rect 63842 222 63894 274
rect 64684 543 64736 552
rect 64684 509 64693 543
rect 64693 509 64727 543
rect 64727 509 64736 543
rect 64684 500 64736 509
rect 65308 667 65360 676
rect 65308 633 65317 667
rect 65317 633 65351 667
rect 65351 633 65360 667
rect 65308 624 65360 633
rect 64902 222 64954 274
rect 65090 222 65142 274
rect 65932 791 65984 800
rect 65932 757 65941 791
rect 65941 757 65975 791
rect 65975 757 65984 791
rect 65932 748 65984 757
rect 66556 419 66608 428
rect 66556 385 66565 419
rect 66565 385 66599 419
rect 66599 385 66608 419
rect 66556 376 66608 385
rect 66150 222 66202 274
rect 66338 222 66390 274
rect 67180 543 67232 552
rect 67180 509 67189 543
rect 67189 509 67223 543
rect 67223 509 67232 543
rect 67180 500 67232 509
rect 67804 667 67856 676
rect 67804 633 67813 667
rect 67813 633 67847 667
rect 67847 633 67856 667
rect 67804 624 67856 633
rect 67398 222 67450 274
rect 67586 222 67638 274
rect 68428 791 68480 800
rect 68428 757 68437 791
rect 68437 757 68471 791
rect 68471 757 68480 791
rect 68428 748 68480 757
rect 69052 419 69104 428
rect 69052 385 69061 419
rect 69061 385 69095 419
rect 69095 385 69104 419
rect 69052 376 69104 385
rect 68646 222 68698 274
rect 68834 222 68886 274
rect 69676 543 69728 552
rect 69676 509 69685 543
rect 69685 509 69719 543
rect 69719 509 69728 543
rect 69676 500 69728 509
rect 70300 667 70352 676
rect 70300 633 70309 667
rect 70309 633 70343 667
rect 70343 633 70352 667
rect 70300 624 70352 633
rect 69894 222 69946 274
rect 70082 222 70134 274
rect 70924 791 70976 800
rect 70924 757 70933 791
rect 70933 757 70967 791
rect 70967 757 70976 791
rect 70924 748 70976 757
rect 71548 419 71600 428
rect 71548 385 71557 419
rect 71557 385 71591 419
rect 71591 385 71600 419
rect 71548 376 71600 385
rect 71142 222 71194 274
rect 71330 222 71382 274
rect 72172 543 72224 552
rect 72172 509 72181 543
rect 72181 509 72215 543
rect 72215 509 72224 543
rect 72172 500 72224 509
rect 72796 667 72848 676
rect 72796 633 72805 667
rect 72805 633 72839 667
rect 72839 633 72848 667
rect 72796 624 72848 633
rect 72390 222 72442 274
rect 72578 222 72630 274
rect 73420 791 73472 800
rect 73420 757 73429 791
rect 73429 757 73463 791
rect 73463 757 73472 791
rect 73420 748 73472 757
rect 74044 419 74096 428
rect 74044 385 74053 419
rect 74053 385 74087 419
rect 74087 385 74096 419
rect 74044 376 74096 385
rect 73638 222 73690 274
rect 73826 222 73878 274
rect 74668 543 74720 552
rect 74668 509 74677 543
rect 74677 509 74711 543
rect 74711 509 74720 543
rect 74668 500 74720 509
rect 75292 667 75344 676
rect 75292 633 75301 667
rect 75301 633 75335 667
rect 75335 633 75344 667
rect 75292 624 75344 633
rect 74886 222 74938 274
rect 75074 222 75126 274
rect 75916 791 75968 800
rect 75916 757 75925 791
rect 75925 757 75959 791
rect 75959 757 75968 791
rect 75916 748 75968 757
rect 76540 419 76592 428
rect 76540 385 76549 419
rect 76549 385 76583 419
rect 76583 385 76592 419
rect 76540 376 76592 385
rect 76134 222 76186 274
rect 76322 222 76374 274
rect 77164 543 77216 552
rect 77164 509 77173 543
rect 77173 509 77207 543
rect 77207 509 77216 543
rect 77164 500 77216 509
rect 77788 667 77840 676
rect 77788 633 77797 667
rect 77797 633 77831 667
rect 77831 633 77840 667
rect 77788 624 77840 633
rect 77382 222 77434 274
rect 77570 222 77622 274
rect 78412 791 78464 800
rect 78412 757 78421 791
rect 78421 757 78455 791
rect 78455 757 78464 791
rect 78412 748 78464 757
rect 79036 419 79088 428
rect 79036 385 79045 419
rect 79045 385 79079 419
rect 79079 385 79088 419
rect 79036 376 79088 385
rect 78630 222 78682 274
rect 78818 222 78870 274
rect 79660 543 79712 552
rect 79660 509 79669 543
rect 79669 509 79703 543
rect 79703 509 79712 543
rect 79660 500 79712 509
rect 80284 667 80336 676
rect 80284 633 80293 667
rect 80293 633 80327 667
rect 80327 633 80336 667
rect 80284 624 80336 633
rect 79878 222 79930 274
rect 80066 222 80118 274
rect 80908 791 80960 800
rect 80908 757 80917 791
rect 80917 757 80951 791
rect 80951 757 80960 791
rect 80908 748 80960 757
rect 81126 222 81178 274
rect 1906 98 1958 150
rect 2038 98 2090 150
rect 3154 98 3206 150
rect 3286 98 3338 150
rect 4402 98 4454 150
rect 4534 98 4586 150
rect 5650 98 5702 150
rect 5782 98 5834 150
rect 6898 98 6950 150
rect 7030 98 7082 150
rect 8146 98 8198 150
rect 8278 98 8330 150
rect 9394 98 9446 150
rect 9526 98 9578 150
rect 10642 98 10694 150
rect 10774 98 10826 150
rect 11890 98 11942 150
rect 12022 98 12074 150
rect 13138 98 13190 150
rect 13270 98 13322 150
rect 14386 98 14438 150
rect 14518 98 14570 150
rect 15634 98 15686 150
rect 15766 98 15818 150
rect 16882 98 16934 150
rect 17014 98 17066 150
rect 18130 98 18182 150
rect 18262 98 18314 150
rect 19378 98 19430 150
rect 19510 98 19562 150
rect 20626 98 20678 150
rect 20758 98 20810 150
rect 21874 98 21926 150
rect 22006 98 22058 150
rect 23122 98 23174 150
rect 23254 98 23306 150
rect 24370 98 24422 150
rect 24502 98 24554 150
rect 25618 98 25670 150
rect 25750 98 25802 150
rect 26866 98 26918 150
rect 26998 98 27050 150
rect 28114 98 28166 150
rect 28246 98 28298 150
rect 29362 98 29414 150
rect 29494 98 29546 150
rect 30610 98 30662 150
rect 30742 98 30794 150
rect 31858 98 31910 150
rect 31990 98 32042 150
rect 33106 98 33158 150
rect 33238 98 33290 150
rect 34354 98 34406 150
rect 34486 98 34538 150
rect 35602 98 35654 150
rect 35734 98 35786 150
rect 36850 98 36902 150
rect 36982 98 37034 150
rect 38098 98 38150 150
rect 38230 98 38282 150
rect 39346 98 39398 150
rect 39478 98 39530 150
rect 40594 98 40646 150
rect 40726 98 40778 150
rect 41842 98 41894 150
rect 41974 98 42026 150
rect 43090 98 43142 150
rect 43222 98 43274 150
rect 44338 98 44390 150
rect 44470 98 44522 150
rect 45586 98 45638 150
rect 45718 98 45770 150
rect 46834 98 46886 150
rect 46966 98 47018 150
rect 48082 98 48134 150
rect 48214 98 48266 150
rect 49330 98 49382 150
rect 49462 98 49514 150
rect 50578 98 50630 150
rect 50710 98 50762 150
rect 51826 98 51878 150
rect 51958 98 52010 150
rect 53074 98 53126 150
rect 53206 98 53258 150
rect 54322 98 54374 150
rect 54454 98 54506 150
rect 55570 98 55622 150
rect 55702 98 55754 150
rect 56818 98 56870 150
rect 56950 98 57002 150
rect 58066 98 58118 150
rect 58198 98 58250 150
rect 59314 98 59366 150
rect 59446 98 59498 150
rect 60562 98 60614 150
rect 60694 98 60746 150
rect 61810 98 61862 150
rect 61942 98 61994 150
rect 63058 98 63110 150
rect 63190 98 63242 150
rect 64306 98 64358 150
rect 64438 98 64490 150
rect 65554 98 65606 150
rect 65686 98 65738 150
rect 66802 98 66854 150
rect 66934 98 66986 150
rect 68050 98 68102 150
rect 68182 98 68234 150
rect 69298 98 69350 150
rect 69430 98 69482 150
rect 70546 98 70598 150
rect 70678 98 70730 150
rect 71794 98 71846 150
rect 71926 98 71978 150
rect 73042 98 73094 150
rect 73174 98 73226 150
rect 74290 98 74342 150
rect 74422 98 74474 150
rect 75538 98 75590 150
rect 75670 98 75722 150
rect 76786 98 76838 150
rect 76918 98 76970 150
rect 78034 98 78086 150
rect 78166 98 78218 150
rect 79282 98 79334 150
rect 79414 98 79466 150
rect 80530 98 80582 150
rect 80662 98 80714 150
<< metal2 >>
rect 3530 802 3586 811
rect 3530 737 3586 746
rect 6026 802 6082 811
rect 6026 737 6082 746
rect 8522 802 8578 811
rect 8522 737 8578 746
rect 11018 802 11074 811
rect 11018 737 11074 746
rect 13514 802 13570 811
rect 13514 737 13570 746
rect 16010 802 16066 811
rect 16010 737 16066 746
rect 18506 802 18562 811
rect 18506 737 18562 746
rect 21002 802 21058 811
rect 21002 737 21058 746
rect 23498 802 23554 811
rect 23498 737 23554 746
rect 25994 802 26050 811
rect 25994 737 26050 746
rect 28490 802 28546 811
rect 28490 737 28546 746
rect 30986 802 31042 811
rect 30986 737 31042 746
rect 33482 802 33538 811
rect 33482 737 33538 746
rect 35978 802 36034 811
rect 35978 737 36034 746
rect 38474 802 38530 811
rect 38474 737 38530 746
rect 40970 802 41026 811
rect 40970 737 41026 746
rect 43466 802 43522 811
rect 43466 737 43522 746
rect 45962 802 46018 811
rect 45962 737 46018 746
rect 48458 802 48514 811
rect 48458 737 48514 746
rect 50954 802 51010 811
rect 50954 737 51010 746
rect 53450 802 53506 811
rect 53450 737 53506 746
rect 55946 802 56002 811
rect 55946 737 56002 746
rect 58442 802 58498 811
rect 58442 737 58498 746
rect 60938 802 60994 811
rect 60938 737 60994 746
rect 63434 802 63490 811
rect 63434 737 63490 746
rect 65930 802 65986 811
rect 65930 737 65986 746
rect 68426 802 68482 811
rect 68426 737 68482 746
rect 70922 802 70978 811
rect 70922 737 70978 746
rect 73418 802 73474 811
rect 73418 737 73474 746
rect 75914 802 75970 811
rect 75914 737 75970 746
rect 78410 802 78466 811
rect 78410 737 78466 746
rect 80906 802 80962 811
rect 80906 737 80962 746
rect 2906 678 2962 687
rect 2906 613 2962 622
rect 5402 678 5458 687
rect 5402 613 5458 622
rect 7898 678 7954 687
rect 7898 613 7954 622
rect 10394 678 10450 687
rect 10394 613 10450 622
rect 12890 678 12946 687
rect 12890 613 12946 622
rect 15386 678 15442 687
rect 15386 613 15442 622
rect 17882 678 17938 687
rect 17882 613 17938 622
rect 20378 678 20434 687
rect 20378 613 20434 622
rect 22874 678 22930 687
rect 22874 613 22930 622
rect 25370 678 25426 687
rect 25370 613 25426 622
rect 27866 678 27922 687
rect 27866 613 27922 622
rect 30362 678 30418 687
rect 30362 613 30418 622
rect 32858 678 32914 687
rect 32858 613 32914 622
rect 35354 678 35410 687
rect 35354 613 35410 622
rect 37850 678 37906 687
rect 37850 613 37906 622
rect 40346 678 40402 687
rect 40346 613 40402 622
rect 42842 678 42898 687
rect 42842 613 42898 622
rect 45338 678 45394 687
rect 45338 613 45394 622
rect 47834 678 47890 687
rect 47834 613 47890 622
rect 50330 678 50386 687
rect 50330 613 50386 622
rect 52826 678 52882 687
rect 52826 613 52882 622
rect 55322 678 55378 687
rect 55322 613 55378 622
rect 57818 678 57874 687
rect 57818 613 57874 622
rect 60314 678 60370 687
rect 60314 613 60370 622
rect 62810 678 62866 687
rect 62810 613 62866 622
rect 65306 678 65362 687
rect 65306 613 65362 622
rect 67802 678 67858 687
rect 67802 613 67858 622
rect 70298 678 70354 687
rect 70298 613 70354 622
rect 72794 678 72850 687
rect 72794 613 72850 622
rect 75290 678 75346 687
rect 75290 613 75346 622
rect 77786 678 77842 687
rect 77786 613 77842 622
rect 80282 678 80338 687
rect 80282 613 80338 622
rect 2282 554 2338 563
rect 2282 489 2338 498
rect 4778 554 4834 563
rect 4778 489 4834 498
rect 7274 554 7330 563
rect 7274 489 7330 498
rect 9770 554 9826 563
rect 9770 489 9826 498
rect 12266 554 12322 563
rect 12266 489 12322 498
rect 14762 554 14818 563
rect 14762 489 14818 498
rect 17258 554 17314 563
rect 17258 489 17314 498
rect 19754 554 19810 563
rect 19754 489 19810 498
rect 22250 554 22306 563
rect 22250 489 22306 498
rect 24746 554 24802 563
rect 24746 489 24802 498
rect 27242 554 27298 563
rect 27242 489 27298 498
rect 29738 554 29794 563
rect 29738 489 29794 498
rect 32234 554 32290 563
rect 32234 489 32290 498
rect 34730 554 34786 563
rect 34730 489 34786 498
rect 37226 554 37282 563
rect 37226 489 37282 498
rect 39722 554 39778 563
rect 39722 489 39778 498
rect 42218 554 42274 563
rect 42218 489 42274 498
rect 44714 554 44770 563
rect 44714 489 44770 498
rect 47210 554 47266 563
rect 47210 489 47266 498
rect 49706 554 49762 563
rect 49706 489 49762 498
rect 52202 554 52258 563
rect 52202 489 52258 498
rect 54698 554 54754 563
rect 54698 489 54754 498
rect 57194 554 57250 563
rect 57194 489 57250 498
rect 59690 554 59746 563
rect 59690 489 59746 498
rect 62186 554 62242 563
rect 62186 489 62242 498
rect 64682 554 64738 563
rect 64682 489 64738 498
rect 67178 554 67234 563
rect 67178 489 67234 498
rect 69674 554 69730 563
rect 69674 489 69730 498
rect 72170 554 72226 563
rect 72170 489 72226 498
rect 74666 554 74722 563
rect 74666 489 74722 498
rect 77162 554 77218 563
rect 77162 489 77218 498
rect 79658 554 79714 563
rect 79658 489 79714 498
rect 1658 430 1714 439
rect 1658 365 1714 374
rect 4154 430 4210 439
rect 4154 365 4210 374
rect 6650 430 6706 439
rect 6650 365 6706 374
rect 9146 430 9202 439
rect 9146 365 9202 374
rect 11642 430 11698 439
rect 11642 365 11698 374
rect 14138 430 14194 439
rect 14138 365 14194 374
rect 16634 430 16690 439
rect 16634 365 16690 374
rect 19130 430 19186 439
rect 19130 365 19186 374
rect 21626 430 21682 439
rect 21626 365 21682 374
rect 24122 430 24178 439
rect 24122 365 24178 374
rect 26618 430 26674 439
rect 26618 365 26674 374
rect 29114 430 29170 439
rect 29114 365 29170 374
rect 31610 430 31666 439
rect 31610 365 31666 374
rect 34106 430 34162 439
rect 34106 365 34162 374
rect 36602 430 36658 439
rect 36602 365 36658 374
rect 39098 430 39154 439
rect 39098 365 39154 374
rect 41594 430 41650 439
rect 41594 365 41650 374
rect 44090 430 44146 439
rect 44090 365 44146 374
rect 46586 430 46642 439
rect 46586 365 46642 374
rect 49082 430 49138 439
rect 49082 365 49138 374
rect 51578 430 51634 439
rect 51578 365 51634 374
rect 54074 430 54130 439
rect 54074 365 54130 374
rect 56570 430 56626 439
rect 56570 365 56626 374
rect 59066 430 59122 439
rect 59066 365 59122 374
rect 61562 430 61618 439
rect 61562 365 61618 374
rect 64058 430 64114 439
rect 64058 365 64114 374
rect 66554 430 66610 439
rect 66554 365 66610 374
rect 69050 430 69106 439
rect 69050 365 69106 374
rect 71546 430 71602 439
rect 71546 365 71602 374
rect 74042 430 74098 439
rect 74042 365 74098 374
rect 76538 430 76594 439
rect 76538 365 76594 374
rect 79034 430 79090 439
rect 79034 365 79090 374
rect 1440 276 1496 285
rect 1440 211 1496 220
rect 2500 276 2556 285
rect 2500 211 2556 220
rect 2688 276 2744 285
rect 2688 211 2744 220
rect 3748 276 3804 285
rect 3748 211 3804 220
rect 3936 276 3992 285
rect 3936 211 3992 220
rect 4996 276 5052 285
rect 4996 211 5052 220
rect 5184 276 5240 285
rect 5184 211 5240 220
rect 6244 276 6300 285
rect 6244 211 6300 220
rect 6432 276 6488 285
rect 6432 211 6488 220
rect 7492 276 7548 285
rect 7492 211 7548 220
rect 7680 276 7736 285
rect 7680 211 7736 220
rect 8740 276 8796 285
rect 8740 211 8796 220
rect 8928 276 8984 285
rect 8928 211 8984 220
rect 9988 276 10044 285
rect 9988 211 10044 220
rect 10176 276 10232 285
rect 10176 211 10232 220
rect 11236 276 11292 285
rect 11236 211 11292 220
rect 11424 276 11480 285
rect 11424 211 11480 220
rect 12484 276 12540 285
rect 12484 211 12540 220
rect 12672 276 12728 285
rect 12672 211 12728 220
rect 13732 276 13788 285
rect 13732 211 13788 220
rect 13920 276 13976 285
rect 13920 211 13976 220
rect 14980 276 15036 285
rect 14980 211 15036 220
rect 15168 276 15224 285
rect 15168 211 15224 220
rect 16228 276 16284 285
rect 16228 211 16284 220
rect 16416 276 16472 285
rect 16416 211 16472 220
rect 17476 276 17532 285
rect 17476 211 17532 220
rect 17664 276 17720 285
rect 17664 211 17720 220
rect 18724 276 18780 285
rect 18724 211 18780 220
rect 18912 276 18968 285
rect 18912 211 18968 220
rect 19972 276 20028 285
rect 19972 211 20028 220
rect 20160 276 20216 285
rect 20160 211 20216 220
rect 21220 276 21276 285
rect 21220 211 21276 220
rect 21408 276 21464 285
rect 21408 211 21464 220
rect 22468 276 22524 285
rect 22468 211 22524 220
rect 22656 276 22712 285
rect 22656 211 22712 220
rect 23716 276 23772 285
rect 23716 211 23772 220
rect 23904 276 23960 285
rect 23904 211 23960 220
rect 24964 276 25020 285
rect 24964 211 25020 220
rect 25152 276 25208 285
rect 25152 211 25208 220
rect 26212 276 26268 285
rect 26212 211 26268 220
rect 26400 276 26456 285
rect 26400 211 26456 220
rect 27460 276 27516 285
rect 27460 211 27516 220
rect 27648 276 27704 285
rect 27648 211 27704 220
rect 28708 276 28764 285
rect 28708 211 28764 220
rect 28896 276 28952 285
rect 28896 211 28952 220
rect 29956 276 30012 285
rect 29956 211 30012 220
rect 30144 276 30200 285
rect 30144 211 30200 220
rect 31204 276 31260 285
rect 31204 211 31260 220
rect 31392 276 31448 285
rect 31392 211 31448 220
rect 32452 276 32508 285
rect 32452 211 32508 220
rect 32640 276 32696 285
rect 32640 211 32696 220
rect 33700 276 33756 285
rect 33700 211 33756 220
rect 33888 276 33944 285
rect 33888 211 33944 220
rect 34948 276 35004 285
rect 34948 211 35004 220
rect 35136 276 35192 285
rect 35136 211 35192 220
rect 36196 276 36252 285
rect 36196 211 36252 220
rect 36384 276 36440 285
rect 36384 211 36440 220
rect 37444 276 37500 285
rect 37444 211 37500 220
rect 37632 276 37688 285
rect 37632 211 37688 220
rect 38692 276 38748 285
rect 38692 211 38748 220
rect 38880 276 38936 285
rect 38880 211 38936 220
rect 39940 276 39996 285
rect 39940 211 39996 220
rect 40128 276 40184 285
rect 40128 211 40184 220
rect 41188 276 41244 285
rect 41188 211 41244 220
rect 41376 276 41432 285
rect 41376 211 41432 220
rect 42436 276 42492 285
rect 42436 211 42492 220
rect 42624 276 42680 285
rect 42624 211 42680 220
rect 43684 276 43740 285
rect 43684 211 43740 220
rect 43872 276 43928 285
rect 43872 211 43928 220
rect 44932 276 44988 285
rect 44932 211 44988 220
rect 45120 276 45176 285
rect 45120 211 45176 220
rect 46180 276 46236 285
rect 46180 211 46236 220
rect 46368 276 46424 285
rect 46368 211 46424 220
rect 47428 276 47484 285
rect 47428 211 47484 220
rect 47616 276 47672 285
rect 47616 211 47672 220
rect 48676 276 48732 285
rect 48676 211 48732 220
rect 48864 276 48920 285
rect 48864 211 48920 220
rect 49924 276 49980 285
rect 49924 211 49980 220
rect 50112 276 50168 285
rect 50112 211 50168 220
rect 51172 276 51228 285
rect 51172 211 51228 220
rect 51360 276 51416 285
rect 51360 211 51416 220
rect 52420 276 52476 285
rect 52420 211 52476 220
rect 52608 276 52664 285
rect 52608 211 52664 220
rect 53668 276 53724 285
rect 53668 211 53724 220
rect 53856 276 53912 285
rect 53856 211 53912 220
rect 54916 276 54972 285
rect 54916 211 54972 220
rect 55104 276 55160 285
rect 55104 211 55160 220
rect 56164 276 56220 285
rect 56164 211 56220 220
rect 56352 276 56408 285
rect 56352 211 56408 220
rect 57412 276 57468 285
rect 57412 211 57468 220
rect 57600 276 57656 285
rect 57600 211 57656 220
rect 58660 276 58716 285
rect 58660 211 58716 220
rect 58848 276 58904 285
rect 58848 211 58904 220
rect 59908 276 59964 285
rect 59908 211 59964 220
rect 60096 276 60152 285
rect 60096 211 60152 220
rect 61156 276 61212 285
rect 61156 211 61212 220
rect 61344 276 61400 285
rect 61344 211 61400 220
rect 62404 276 62460 285
rect 62404 211 62460 220
rect 62592 276 62648 285
rect 62592 211 62648 220
rect 63652 276 63708 285
rect 63652 211 63708 220
rect 63840 276 63896 285
rect 63840 211 63896 220
rect 64900 276 64956 285
rect 64900 211 64956 220
rect 65088 276 65144 285
rect 65088 211 65144 220
rect 66148 276 66204 285
rect 66148 211 66204 220
rect 66336 276 66392 285
rect 66336 211 66392 220
rect 67396 276 67452 285
rect 67396 211 67452 220
rect 67584 276 67640 285
rect 67584 211 67640 220
rect 68644 276 68700 285
rect 68644 211 68700 220
rect 68832 276 68888 285
rect 68832 211 68888 220
rect 69892 276 69948 285
rect 69892 211 69948 220
rect 70080 276 70136 285
rect 70080 211 70136 220
rect 71140 276 71196 285
rect 71140 211 71196 220
rect 71328 276 71384 285
rect 71328 211 71384 220
rect 72388 276 72444 285
rect 72388 211 72444 220
rect 72576 276 72632 285
rect 72576 211 72632 220
rect 73636 276 73692 285
rect 73636 211 73692 220
rect 73824 276 73880 285
rect 73824 211 73880 220
rect 74884 276 74940 285
rect 74884 211 74940 220
rect 75072 276 75128 285
rect 75072 211 75128 220
rect 76132 276 76188 285
rect 76132 211 76188 220
rect 76320 276 76376 285
rect 76320 211 76376 220
rect 77380 276 77436 285
rect 77380 211 77436 220
rect 77568 276 77624 285
rect 77568 211 77624 220
rect 78628 276 78684 285
rect 78628 211 78684 220
rect 78816 276 78872 285
rect 78816 211 78872 220
rect 79876 276 79932 285
rect 79876 211 79932 220
rect 80064 276 80120 285
rect 80064 211 80120 220
rect 81124 276 81180 285
rect 81124 211 81180 220
rect 1904 152 1960 161
rect 1904 87 1960 96
rect 2036 152 2092 161
rect 2036 87 2092 96
rect 3152 152 3208 161
rect 3152 87 3208 96
rect 3284 152 3340 161
rect 3284 87 3340 96
rect 4400 152 4456 161
rect 4400 87 4456 96
rect 4532 152 4588 161
rect 4532 87 4588 96
rect 5648 152 5704 161
rect 5648 87 5704 96
rect 5780 152 5836 161
rect 5780 87 5836 96
rect 6896 152 6952 161
rect 6896 87 6952 96
rect 7028 152 7084 161
rect 7028 87 7084 96
rect 8144 152 8200 161
rect 8144 87 8200 96
rect 8276 152 8332 161
rect 8276 87 8332 96
rect 9392 152 9448 161
rect 9392 87 9448 96
rect 9524 152 9580 161
rect 9524 87 9580 96
rect 10640 152 10696 161
rect 10640 87 10696 96
rect 10772 152 10828 161
rect 10772 87 10828 96
rect 11888 152 11944 161
rect 11888 87 11944 96
rect 12020 152 12076 161
rect 12020 87 12076 96
rect 13136 152 13192 161
rect 13136 87 13192 96
rect 13268 152 13324 161
rect 13268 87 13324 96
rect 14384 152 14440 161
rect 14384 87 14440 96
rect 14516 152 14572 161
rect 14516 87 14572 96
rect 15632 152 15688 161
rect 15632 87 15688 96
rect 15764 152 15820 161
rect 15764 87 15820 96
rect 16880 152 16936 161
rect 16880 87 16936 96
rect 17012 152 17068 161
rect 17012 87 17068 96
rect 18128 152 18184 161
rect 18128 87 18184 96
rect 18260 152 18316 161
rect 18260 87 18316 96
rect 19376 152 19432 161
rect 19376 87 19432 96
rect 19508 152 19564 161
rect 19508 87 19564 96
rect 20624 152 20680 161
rect 20624 87 20680 96
rect 20756 152 20812 161
rect 20756 87 20812 96
rect 21872 152 21928 161
rect 21872 87 21928 96
rect 22004 152 22060 161
rect 22004 87 22060 96
rect 23120 152 23176 161
rect 23120 87 23176 96
rect 23252 152 23308 161
rect 23252 87 23308 96
rect 24368 152 24424 161
rect 24368 87 24424 96
rect 24500 152 24556 161
rect 24500 87 24556 96
rect 25616 152 25672 161
rect 25616 87 25672 96
rect 25748 152 25804 161
rect 25748 87 25804 96
rect 26864 152 26920 161
rect 26864 87 26920 96
rect 26996 152 27052 161
rect 26996 87 27052 96
rect 28112 152 28168 161
rect 28112 87 28168 96
rect 28244 152 28300 161
rect 28244 87 28300 96
rect 29360 152 29416 161
rect 29360 87 29416 96
rect 29492 152 29548 161
rect 29492 87 29548 96
rect 30608 152 30664 161
rect 30608 87 30664 96
rect 30740 152 30796 161
rect 30740 87 30796 96
rect 31856 152 31912 161
rect 31856 87 31912 96
rect 31988 152 32044 161
rect 31988 87 32044 96
rect 33104 152 33160 161
rect 33104 87 33160 96
rect 33236 152 33292 161
rect 33236 87 33292 96
rect 34352 152 34408 161
rect 34352 87 34408 96
rect 34484 152 34540 161
rect 34484 87 34540 96
rect 35600 152 35656 161
rect 35600 87 35656 96
rect 35732 152 35788 161
rect 35732 87 35788 96
rect 36848 152 36904 161
rect 36848 87 36904 96
rect 36980 152 37036 161
rect 36980 87 37036 96
rect 38096 152 38152 161
rect 38096 87 38152 96
rect 38228 152 38284 161
rect 38228 87 38284 96
rect 39344 152 39400 161
rect 39344 87 39400 96
rect 39476 152 39532 161
rect 39476 87 39532 96
rect 40592 152 40648 161
rect 40592 87 40648 96
rect 40724 152 40780 161
rect 40724 87 40780 96
rect 41840 152 41896 161
rect 41840 87 41896 96
rect 41972 152 42028 161
rect 41972 87 42028 96
rect 43088 152 43144 161
rect 43088 87 43144 96
rect 43220 152 43276 161
rect 43220 87 43276 96
rect 44336 152 44392 161
rect 44336 87 44392 96
rect 44468 152 44524 161
rect 44468 87 44524 96
rect 45584 152 45640 161
rect 45584 87 45640 96
rect 45716 152 45772 161
rect 45716 87 45772 96
rect 46832 152 46888 161
rect 46832 87 46888 96
rect 46964 152 47020 161
rect 46964 87 47020 96
rect 48080 152 48136 161
rect 48080 87 48136 96
rect 48212 152 48268 161
rect 48212 87 48268 96
rect 49328 152 49384 161
rect 49328 87 49384 96
rect 49460 152 49516 161
rect 49460 87 49516 96
rect 50576 152 50632 161
rect 50576 87 50632 96
rect 50708 152 50764 161
rect 50708 87 50764 96
rect 51824 152 51880 161
rect 51824 87 51880 96
rect 51956 152 52012 161
rect 51956 87 52012 96
rect 53072 152 53128 161
rect 53072 87 53128 96
rect 53204 152 53260 161
rect 53204 87 53260 96
rect 54320 152 54376 161
rect 54320 87 54376 96
rect 54452 152 54508 161
rect 54452 87 54508 96
rect 55568 152 55624 161
rect 55568 87 55624 96
rect 55700 152 55756 161
rect 55700 87 55756 96
rect 56816 152 56872 161
rect 56816 87 56872 96
rect 56948 152 57004 161
rect 56948 87 57004 96
rect 58064 152 58120 161
rect 58064 87 58120 96
rect 58196 152 58252 161
rect 58196 87 58252 96
rect 59312 152 59368 161
rect 59312 87 59368 96
rect 59444 152 59500 161
rect 59444 87 59500 96
rect 60560 152 60616 161
rect 60560 87 60616 96
rect 60692 152 60748 161
rect 60692 87 60748 96
rect 61808 152 61864 161
rect 61808 87 61864 96
rect 61940 152 61996 161
rect 61940 87 61996 96
rect 63056 152 63112 161
rect 63056 87 63112 96
rect 63188 152 63244 161
rect 63188 87 63244 96
rect 64304 152 64360 161
rect 64304 87 64360 96
rect 64436 152 64492 161
rect 64436 87 64492 96
rect 65552 152 65608 161
rect 65552 87 65608 96
rect 65684 152 65740 161
rect 65684 87 65740 96
rect 66800 152 66856 161
rect 66800 87 66856 96
rect 66932 152 66988 161
rect 66932 87 66988 96
rect 68048 152 68104 161
rect 68048 87 68104 96
rect 68180 152 68236 161
rect 68180 87 68236 96
rect 69296 152 69352 161
rect 69296 87 69352 96
rect 69428 152 69484 161
rect 69428 87 69484 96
rect 70544 152 70600 161
rect 70544 87 70600 96
rect 70676 152 70732 161
rect 70676 87 70732 96
rect 71792 152 71848 161
rect 71792 87 71848 96
rect 71924 152 71980 161
rect 71924 87 71980 96
rect 73040 152 73096 161
rect 73040 87 73096 96
rect 73172 152 73228 161
rect 73172 87 73228 96
rect 74288 152 74344 161
rect 74288 87 74344 96
rect 74420 152 74476 161
rect 74420 87 74476 96
rect 75536 152 75592 161
rect 75536 87 75592 96
rect 75668 152 75724 161
rect 75668 87 75724 96
rect 76784 152 76840 161
rect 76784 87 76840 96
rect 76916 152 76972 161
rect 76916 87 76972 96
rect 78032 152 78088 161
rect 78032 87 78088 96
rect 78164 152 78220 161
rect 78164 87 78220 96
rect 79280 152 79336 161
rect 79280 87 79336 96
rect 79412 152 79468 161
rect 79412 87 79468 96
rect 80528 152 80584 161
rect 80528 87 80584 96
rect 80660 152 80716 161
rect 80660 87 80716 96
<< via2 >>
rect 3530 800 3586 802
rect 3530 748 3532 800
rect 3532 748 3584 800
rect 3584 748 3586 800
rect 3530 746 3586 748
rect 6026 800 6082 802
rect 6026 748 6028 800
rect 6028 748 6080 800
rect 6080 748 6082 800
rect 6026 746 6082 748
rect 8522 800 8578 802
rect 8522 748 8524 800
rect 8524 748 8576 800
rect 8576 748 8578 800
rect 8522 746 8578 748
rect 11018 800 11074 802
rect 11018 748 11020 800
rect 11020 748 11072 800
rect 11072 748 11074 800
rect 11018 746 11074 748
rect 13514 800 13570 802
rect 13514 748 13516 800
rect 13516 748 13568 800
rect 13568 748 13570 800
rect 13514 746 13570 748
rect 16010 800 16066 802
rect 16010 748 16012 800
rect 16012 748 16064 800
rect 16064 748 16066 800
rect 16010 746 16066 748
rect 18506 800 18562 802
rect 18506 748 18508 800
rect 18508 748 18560 800
rect 18560 748 18562 800
rect 18506 746 18562 748
rect 21002 800 21058 802
rect 21002 748 21004 800
rect 21004 748 21056 800
rect 21056 748 21058 800
rect 21002 746 21058 748
rect 23498 800 23554 802
rect 23498 748 23500 800
rect 23500 748 23552 800
rect 23552 748 23554 800
rect 23498 746 23554 748
rect 25994 800 26050 802
rect 25994 748 25996 800
rect 25996 748 26048 800
rect 26048 748 26050 800
rect 25994 746 26050 748
rect 28490 800 28546 802
rect 28490 748 28492 800
rect 28492 748 28544 800
rect 28544 748 28546 800
rect 28490 746 28546 748
rect 30986 800 31042 802
rect 30986 748 30988 800
rect 30988 748 31040 800
rect 31040 748 31042 800
rect 30986 746 31042 748
rect 33482 800 33538 802
rect 33482 748 33484 800
rect 33484 748 33536 800
rect 33536 748 33538 800
rect 33482 746 33538 748
rect 35978 800 36034 802
rect 35978 748 35980 800
rect 35980 748 36032 800
rect 36032 748 36034 800
rect 35978 746 36034 748
rect 38474 800 38530 802
rect 38474 748 38476 800
rect 38476 748 38528 800
rect 38528 748 38530 800
rect 38474 746 38530 748
rect 40970 800 41026 802
rect 40970 748 40972 800
rect 40972 748 41024 800
rect 41024 748 41026 800
rect 40970 746 41026 748
rect 43466 800 43522 802
rect 43466 748 43468 800
rect 43468 748 43520 800
rect 43520 748 43522 800
rect 43466 746 43522 748
rect 45962 800 46018 802
rect 45962 748 45964 800
rect 45964 748 46016 800
rect 46016 748 46018 800
rect 45962 746 46018 748
rect 48458 800 48514 802
rect 48458 748 48460 800
rect 48460 748 48512 800
rect 48512 748 48514 800
rect 48458 746 48514 748
rect 50954 800 51010 802
rect 50954 748 50956 800
rect 50956 748 51008 800
rect 51008 748 51010 800
rect 50954 746 51010 748
rect 53450 800 53506 802
rect 53450 748 53452 800
rect 53452 748 53504 800
rect 53504 748 53506 800
rect 53450 746 53506 748
rect 55946 800 56002 802
rect 55946 748 55948 800
rect 55948 748 56000 800
rect 56000 748 56002 800
rect 55946 746 56002 748
rect 58442 800 58498 802
rect 58442 748 58444 800
rect 58444 748 58496 800
rect 58496 748 58498 800
rect 58442 746 58498 748
rect 60938 800 60994 802
rect 60938 748 60940 800
rect 60940 748 60992 800
rect 60992 748 60994 800
rect 60938 746 60994 748
rect 63434 800 63490 802
rect 63434 748 63436 800
rect 63436 748 63488 800
rect 63488 748 63490 800
rect 63434 746 63490 748
rect 65930 800 65986 802
rect 65930 748 65932 800
rect 65932 748 65984 800
rect 65984 748 65986 800
rect 65930 746 65986 748
rect 68426 800 68482 802
rect 68426 748 68428 800
rect 68428 748 68480 800
rect 68480 748 68482 800
rect 68426 746 68482 748
rect 70922 800 70978 802
rect 70922 748 70924 800
rect 70924 748 70976 800
rect 70976 748 70978 800
rect 70922 746 70978 748
rect 73418 800 73474 802
rect 73418 748 73420 800
rect 73420 748 73472 800
rect 73472 748 73474 800
rect 73418 746 73474 748
rect 75914 800 75970 802
rect 75914 748 75916 800
rect 75916 748 75968 800
rect 75968 748 75970 800
rect 75914 746 75970 748
rect 78410 800 78466 802
rect 78410 748 78412 800
rect 78412 748 78464 800
rect 78464 748 78466 800
rect 78410 746 78466 748
rect 80906 800 80962 802
rect 80906 748 80908 800
rect 80908 748 80960 800
rect 80960 748 80962 800
rect 80906 746 80962 748
rect 2906 676 2962 678
rect 2906 624 2908 676
rect 2908 624 2960 676
rect 2960 624 2962 676
rect 2906 622 2962 624
rect 5402 676 5458 678
rect 5402 624 5404 676
rect 5404 624 5456 676
rect 5456 624 5458 676
rect 5402 622 5458 624
rect 7898 676 7954 678
rect 7898 624 7900 676
rect 7900 624 7952 676
rect 7952 624 7954 676
rect 7898 622 7954 624
rect 10394 676 10450 678
rect 10394 624 10396 676
rect 10396 624 10448 676
rect 10448 624 10450 676
rect 10394 622 10450 624
rect 12890 676 12946 678
rect 12890 624 12892 676
rect 12892 624 12944 676
rect 12944 624 12946 676
rect 12890 622 12946 624
rect 15386 676 15442 678
rect 15386 624 15388 676
rect 15388 624 15440 676
rect 15440 624 15442 676
rect 15386 622 15442 624
rect 17882 676 17938 678
rect 17882 624 17884 676
rect 17884 624 17936 676
rect 17936 624 17938 676
rect 17882 622 17938 624
rect 20378 676 20434 678
rect 20378 624 20380 676
rect 20380 624 20432 676
rect 20432 624 20434 676
rect 20378 622 20434 624
rect 22874 676 22930 678
rect 22874 624 22876 676
rect 22876 624 22928 676
rect 22928 624 22930 676
rect 22874 622 22930 624
rect 25370 676 25426 678
rect 25370 624 25372 676
rect 25372 624 25424 676
rect 25424 624 25426 676
rect 25370 622 25426 624
rect 27866 676 27922 678
rect 27866 624 27868 676
rect 27868 624 27920 676
rect 27920 624 27922 676
rect 27866 622 27922 624
rect 30362 676 30418 678
rect 30362 624 30364 676
rect 30364 624 30416 676
rect 30416 624 30418 676
rect 30362 622 30418 624
rect 32858 676 32914 678
rect 32858 624 32860 676
rect 32860 624 32912 676
rect 32912 624 32914 676
rect 32858 622 32914 624
rect 35354 676 35410 678
rect 35354 624 35356 676
rect 35356 624 35408 676
rect 35408 624 35410 676
rect 35354 622 35410 624
rect 37850 676 37906 678
rect 37850 624 37852 676
rect 37852 624 37904 676
rect 37904 624 37906 676
rect 37850 622 37906 624
rect 40346 676 40402 678
rect 40346 624 40348 676
rect 40348 624 40400 676
rect 40400 624 40402 676
rect 40346 622 40402 624
rect 42842 676 42898 678
rect 42842 624 42844 676
rect 42844 624 42896 676
rect 42896 624 42898 676
rect 42842 622 42898 624
rect 45338 676 45394 678
rect 45338 624 45340 676
rect 45340 624 45392 676
rect 45392 624 45394 676
rect 45338 622 45394 624
rect 47834 676 47890 678
rect 47834 624 47836 676
rect 47836 624 47888 676
rect 47888 624 47890 676
rect 47834 622 47890 624
rect 50330 676 50386 678
rect 50330 624 50332 676
rect 50332 624 50384 676
rect 50384 624 50386 676
rect 50330 622 50386 624
rect 52826 676 52882 678
rect 52826 624 52828 676
rect 52828 624 52880 676
rect 52880 624 52882 676
rect 52826 622 52882 624
rect 55322 676 55378 678
rect 55322 624 55324 676
rect 55324 624 55376 676
rect 55376 624 55378 676
rect 55322 622 55378 624
rect 57818 676 57874 678
rect 57818 624 57820 676
rect 57820 624 57872 676
rect 57872 624 57874 676
rect 57818 622 57874 624
rect 60314 676 60370 678
rect 60314 624 60316 676
rect 60316 624 60368 676
rect 60368 624 60370 676
rect 60314 622 60370 624
rect 62810 676 62866 678
rect 62810 624 62812 676
rect 62812 624 62864 676
rect 62864 624 62866 676
rect 62810 622 62866 624
rect 65306 676 65362 678
rect 65306 624 65308 676
rect 65308 624 65360 676
rect 65360 624 65362 676
rect 65306 622 65362 624
rect 67802 676 67858 678
rect 67802 624 67804 676
rect 67804 624 67856 676
rect 67856 624 67858 676
rect 67802 622 67858 624
rect 70298 676 70354 678
rect 70298 624 70300 676
rect 70300 624 70352 676
rect 70352 624 70354 676
rect 70298 622 70354 624
rect 72794 676 72850 678
rect 72794 624 72796 676
rect 72796 624 72848 676
rect 72848 624 72850 676
rect 72794 622 72850 624
rect 75290 676 75346 678
rect 75290 624 75292 676
rect 75292 624 75344 676
rect 75344 624 75346 676
rect 75290 622 75346 624
rect 77786 676 77842 678
rect 77786 624 77788 676
rect 77788 624 77840 676
rect 77840 624 77842 676
rect 77786 622 77842 624
rect 80282 676 80338 678
rect 80282 624 80284 676
rect 80284 624 80336 676
rect 80336 624 80338 676
rect 80282 622 80338 624
rect 2282 552 2338 554
rect 2282 500 2284 552
rect 2284 500 2336 552
rect 2336 500 2338 552
rect 2282 498 2338 500
rect 4778 552 4834 554
rect 4778 500 4780 552
rect 4780 500 4832 552
rect 4832 500 4834 552
rect 4778 498 4834 500
rect 7274 552 7330 554
rect 7274 500 7276 552
rect 7276 500 7328 552
rect 7328 500 7330 552
rect 7274 498 7330 500
rect 9770 552 9826 554
rect 9770 500 9772 552
rect 9772 500 9824 552
rect 9824 500 9826 552
rect 9770 498 9826 500
rect 12266 552 12322 554
rect 12266 500 12268 552
rect 12268 500 12320 552
rect 12320 500 12322 552
rect 12266 498 12322 500
rect 14762 552 14818 554
rect 14762 500 14764 552
rect 14764 500 14816 552
rect 14816 500 14818 552
rect 14762 498 14818 500
rect 17258 552 17314 554
rect 17258 500 17260 552
rect 17260 500 17312 552
rect 17312 500 17314 552
rect 17258 498 17314 500
rect 19754 552 19810 554
rect 19754 500 19756 552
rect 19756 500 19808 552
rect 19808 500 19810 552
rect 19754 498 19810 500
rect 22250 552 22306 554
rect 22250 500 22252 552
rect 22252 500 22304 552
rect 22304 500 22306 552
rect 22250 498 22306 500
rect 24746 552 24802 554
rect 24746 500 24748 552
rect 24748 500 24800 552
rect 24800 500 24802 552
rect 24746 498 24802 500
rect 27242 552 27298 554
rect 27242 500 27244 552
rect 27244 500 27296 552
rect 27296 500 27298 552
rect 27242 498 27298 500
rect 29738 552 29794 554
rect 29738 500 29740 552
rect 29740 500 29792 552
rect 29792 500 29794 552
rect 29738 498 29794 500
rect 32234 552 32290 554
rect 32234 500 32236 552
rect 32236 500 32288 552
rect 32288 500 32290 552
rect 32234 498 32290 500
rect 34730 552 34786 554
rect 34730 500 34732 552
rect 34732 500 34784 552
rect 34784 500 34786 552
rect 34730 498 34786 500
rect 37226 552 37282 554
rect 37226 500 37228 552
rect 37228 500 37280 552
rect 37280 500 37282 552
rect 37226 498 37282 500
rect 39722 552 39778 554
rect 39722 500 39724 552
rect 39724 500 39776 552
rect 39776 500 39778 552
rect 39722 498 39778 500
rect 42218 552 42274 554
rect 42218 500 42220 552
rect 42220 500 42272 552
rect 42272 500 42274 552
rect 42218 498 42274 500
rect 44714 552 44770 554
rect 44714 500 44716 552
rect 44716 500 44768 552
rect 44768 500 44770 552
rect 44714 498 44770 500
rect 47210 552 47266 554
rect 47210 500 47212 552
rect 47212 500 47264 552
rect 47264 500 47266 552
rect 47210 498 47266 500
rect 49706 552 49762 554
rect 49706 500 49708 552
rect 49708 500 49760 552
rect 49760 500 49762 552
rect 49706 498 49762 500
rect 52202 552 52258 554
rect 52202 500 52204 552
rect 52204 500 52256 552
rect 52256 500 52258 552
rect 52202 498 52258 500
rect 54698 552 54754 554
rect 54698 500 54700 552
rect 54700 500 54752 552
rect 54752 500 54754 552
rect 54698 498 54754 500
rect 57194 552 57250 554
rect 57194 500 57196 552
rect 57196 500 57248 552
rect 57248 500 57250 552
rect 57194 498 57250 500
rect 59690 552 59746 554
rect 59690 500 59692 552
rect 59692 500 59744 552
rect 59744 500 59746 552
rect 59690 498 59746 500
rect 62186 552 62242 554
rect 62186 500 62188 552
rect 62188 500 62240 552
rect 62240 500 62242 552
rect 62186 498 62242 500
rect 64682 552 64738 554
rect 64682 500 64684 552
rect 64684 500 64736 552
rect 64736 500 64738 552
rect 64682 498 64738 500
rect 67178 552 67234 554
rect 67178 500 67180 552
rect 67180 500 67232 552
rect 67232 500 67234 552
rect 67178 498 67234 500
rect 69674 552 69730 554
rect 69674 500 69676 552
rect 69676 500 69728 552
rect 69728 500 69730 552
rect 69674 498 69730 500
rect 72170 552 72226 554
rect 72170 500 72172 552
rect 72172 500 72224 552
rect 72224 500 72226 552
rect 72170 498 72226 500
rect 74666 552 74722 554
rect 74666 500 74668 552
rect 74668 500 74720 552
rect 74720 500 74722 552
rect 74666 498 74722 500
rect 77162 552 77218 554
rect 77162 500 77164 552
rect 77164 500 77216 552
rect 77216 500 77218 552
rect 77162 498 77218 500
rect 79658 552 79714 554
rect 79658 500 79660 552
rect 79660 500 79712 552
rect 79712 500 79714 552
rect 79658 498 79714 500
rect 1658 428 1714 430
rect 1658 376 1660 428
rect 1660 376 1712 428
rect 1712 376 1714 428
rect 1658 374 1714 376
rect 4154 428 4210 430
rect 4154 376 4156 428
rect 4156 376 4208 428
rect 4208 376 4210 428
rect 4154 374 4210 376
rect 6650 428 6706 430
rect 6650 376 6652 428
rect 6652 376 6704 428
rect 6704 376 6706 428
rect 6650 374 6706 376
rect 9146 428 9202 430
rect 9146 376 9148 428
rect 9148 376 9200 428
rect 9200 376 9202 428
rect 9146 374 9202 376
rect 11642 428 11698 430
rect 11642 376 11644 428
rect 11644 376 11696 428
rect 11696 376 11698 428
rect 11642 374 11698 376
rect 14138 428 14194 430
rect 14138 376 14140 428
rect 14140 376 14192 428
rect 14192 376 14194 428
rect 14138 374 14194 376
rect 16634 428 16690 430
rect 16634 376 16636 428
rect 16636 376 16688 428
rect 16688 376 16690 428
rect 16634 374 16690 376
rect 19130 428 19186 430
rect 19130 376 19132 428
rect 19132 376 19184 428
rect 19184 376 19186 428
rect 19130 374 19186 376
rect 21626 428 21682 430
rect 21626 376 21628 428
rect 21628 376 21680 428
rect 21680 376 21682 428
rect 21626 374 21682 376
rect 24122 428 24178 430
rect 24122 376 24124 428
rect 24124 376 24176 428
rect 24176 376 24178 428
rect 24122 374 24178 376
rect 26618 428 26674 430
rect 26618 376 26620 428
rect 26620 376 26672 428
rect 26672 376 26674 428
rect 26618 374 26674 376
rect 29114 428 29170 430
rect 29114 376 29116 428
rect 29116 376 29168 428
rect 29168 376 29170 428
rect 29114 374 29170 376
rect 31610 428 31666 430
rect 31610 376 31612 428
rect 31612 376 31664 428
rect 31664 376 31666 428
rect 31610 374 31666 376
rect 34106 428 34162 430
rect 34106 376 34108 428
rect 34108 376 34160 428
rect 34160 376 34162 428
rect 34106 374 34162 376
rect 36602 428 36658 430
rect 36602 376 36604 428
rect 36604 376 36656 428
rect 36656 376 36658 428
rect 36602 374 36658 376
rect 39098 428 39154 430
rect 39098 376 39100 428
rect 39100 376 39152 428
rect 39152 376 39154 428
rect 39098 374 39154 376
rect 41594 428 41650 430
rect 41594 376 41596 428
rect 41596 376 41648 428
rect 41648 376 41650 428
rect 41594 374 41650 376
rect 44090 428 44146 430
rect 44090 376 44092 428
rect 44092 376 44144 428
rect 44144 376 44146 428
rect 44090 374 44146 376
rect 46586 428 46642 430
rect 46586 376 46588 428
rect 46588 376 46640 428
rect 46640 376 46642 428
rect 46586 374 46642 376
rect 49082 428 49138 430
rect 49082 376 49084 428
rect 49084 376 49136 428
rect 49136 376 49138 428
rect 49082 374 49138 376
rect 51578 428 51634 430
rect 51578 376 51580 428
rect 51580 376 51632 428
rect 51632 376 51634 428
rect 51578 374 51634 376
rect 54074 428 54130 430
rect 54074 376 54076 428
rect 54076 376 54128 428
rect 54128 376 54130 428
rect 54074 374 54130 376
rect 56570 428 56626 430
rect 56570 376 56572 428
rect 56572 376 56624 428
rect 56624 376 56626 428
rect 56570 374 56626 376
rect 59066 428 59122 430
rect 59066 376 59068 428
rect 59068 376 59120 428
rect 59120 376 59122 428
rect 59066 374 59122 376
rect 61562 428 61618 430
rect 61562 376 61564 428
rect 61564 376 61616 428
rect 61616 376 61618 428
rect 61562 374 61618 376
rect 64058 428 64114 430
rect 64058 376 64060 428
rect 64060 376 64112 428
rect 64112 376 64114 428
rect 64058 374 64114 376
rect 66554 428 66610 430
rect 66554 376 66556 428
rect 66556 376 66608 428
rect 66608 376 66610 428
rect 66554 374 66610 376
rect 69050 428 69106 430
rect 69050 376 69052 428
rect 69052 376 69104 428
rect 69104 376 69106 428
rect 69050 374 69106 376
rect 71546 428 71602 430
rect 71546 376 71548 428
rect 71548 376 71600 428
rect 71600 376 71602 428
rect 71546 374 71602 376
rect 74042 428 74098 430
rect 74042 376 74044 428
rect 74044 376 74096 428
rect 74096 376 74098 428
rect 74042 374 74098 376
rect 76538 428 76594 430
rect 76538 376 76540 428
rect 76540 376 76592 428
rect 76592 376 76594 428
rect 76538 374 76594 376
rect 79034 428 79090 430
rect 79034 376 79036 428
rect 79036 376 79088 428
rect 79088 376 79090 428
rect 79034 374 79090 376
rect 1440 274 1496 276
rect 1440 222 1442 274
rect 1442 222 1494 274
rect 1494 222 1496 274
rect 1440 220 1496 222
rect 2500 274 2556 276
rect 2500 222 2502 274
rect 2502 222 2554 274
rect 2554 222 2556 274
rect 2500 220 2556 222
rect 2688 274 2744 276
rect 2688 222 2690 274
rect 2690 222 2742 274
rect 2742 222 2744 274
rect 2688 220 2744 222
rect 3748 274 3804 276
rect 3748 222 3750 274
rect 3750 222 3802 274
rect 3802 222 3804 274
rect 3748 220 3804 222
rect 3936 274 3992 276
rect 3936 222 3938 274
rect 3938 222 3990 274
rect 3990 222 3992 274
rect 3936 220 3992 222
rect 4996 274 5052 276
rect 4996 222 4998 274
rect 4998 222 5050 274
rect 5050 222 5052 274
rect 4996 220 5052 222
rect 5184 274 5240 276
rect 5184 222 5186 274
rect 5186 222 5238 274
rect 5238 222 5240 274
rect 5184 220 5240 222
rect 6244 274 6300 276
rect 6244 222 6246 274
rect 6246 222 6298 274
rect 6298 222 6300 274
rect 6244 220 6300 222
rect 6432 274 6488 276
rect 6432 222 6434 274
rect 6434 222 6486 274
rect 6486 222 6488 274
rect 6432 220 6488 222
rect 7492 274 7548 276
rect 7492 222 7494 274
rect 7494 222 7546 274
rect 7546 222 7548 274
rect 7492 220 7548 222
rect 7680 274 7736 276
rect 7680 222 7682 274
rect 7682 222 7734 274
rect 7734 222 7736 274
rect 7680 220 7736 222
rect 8740 274 8796 276
rect 8740 222 8742 274
rect 8742 222 8794 274
rect 8794 222 8796 274
rect 8740 220 8796 222
rect 8928 274 8984 276
rect 8928 222 8930 274
rect 8930 222 8982 274
rect 8982 222 8984 274
rect 8928 220 8984 222
rect 9988 274 10044 276
rect 9988 222 9990 274
rect 9990 222 10042 274
rect 10042 222 10044 274
rect 9988 220 10044 222
rect 10176 274 10232 276
rect 10176 222 10178 274
rect 10178 222 10230 274
rect 10230 222 10232 274
rect 10176 220 10232 222
rect 11236 274 11292 276
rect 11236 222 11238 274
rect 11238 222 11290 274
rect 11290 222 11292 274
rect 11236 220 11292 222
rect 11424 274 11480 276
rect 11424 222 11426 274
rect 11426 222 11478 274
rect 11478 222 11480 274
rect 11424 220 11480 222
rect 12484 274 12540 276
rect 12484 222 12486 274
rect 12486 222 12538 274
rect 12538 222 12540 274
rect 12484 220 12540 222
rect 12672 274 12728 276
rect 12672 222 12674 274
rect 12674 222 12726 274
rect 12726 222 12728 274
rect 12672 220 12728 222
rect 13732 274 13788 276
rect 13732 222 13734 274
rect 13734 222 13786 274
rect 13786 222 13788 274
rect 13732 220 13788 222
rect 13920 274 13976 276
rect 13920 222 13922 274
rect 13922 222 13974 274
rect 13974 222 13976 274
rect 13920 220 13976 222
rect 14980 274 15036 276
rect 14980 222 14982 274
rect 14982 222 15034 274
rect 15034 222 15036 274
rect 14980 220 15036 222
rect 15168 274 15224 276
rect 15168 222 15170 274
rect 15170 222 15222 274
rect 15222 222 15224 274
rect 15168 220 15224 222
rect 16228 274 16284 276
rect 16228 222 16230 274
rect 16230 222 16282 274
rect 16282 222 16284 274
rect 16228 220 16284 222
rect 16416 274 16472 276
rect 16416 222 16418 274
rect 16418 222 16470 274
rect 16470 222 16472 274
rect 16416 220 16472 222
rect 17476 274 17532 276
rect 17476 222 17478 274
rect 17478 222 17530 274
rect 17530 222 17532 274
rect 17476 220 17532 222
rect 17664 274 17720 276
rect 17664 222 17666 274
rect 17666 222 17718 274
rect 17718 222 17720 274
rect 17664 220 17720 222
rect 18724 274 18780 276
rect 18724 222 18726 274
rect 18726 222 18778 274
rect 18778 222 18780 274
rect 18724 220 18780 222
rect 18912 274 18968 276
rect 18912 222 18914 274
rect 18914 222 18966 274
rect 18966 222 18968 274
rect 18912 220 18968 222
rect 19972 274 20028 276
rect 19972 222 19974 274
rect 19974 222 20026 274
rect 20026 222 20028 274
rect 19972 220 20028 222
rect 20160 274 20216 276
rect 20160 222 20162 274
rect 20162 222 20214 274
rect 20214 222 20216 274
rect 20160 220 20216 222
rect 21220 274 21276 276
rect 21220 222 21222 274
rect 21222 222 21274 274
rect 21274 222 21276 274
rect 21220 220 21276 222
rect 21408 274 21464 276
rect 21408 222 21410 274
rect 21410 222 21462 274
rect 21462 222 21464 274
rect 21408 220 21464 222
rect 22468 274 22524 276
rect 22468 222 22470 274
rect 22470 222 22522 274
rect 22522 222 22524 274
rect 22468 220 22524 222
rect 22656 274 22712 276
rect 22656 222 22658 274
rect 22658 222 22710 274
rect 22710 222 22712 274
rect 22656 220 22712 222
rect 23716 274 23772 276
rect 23716 222 23718 274
rect 23718 222 23770 274
rect 23770 222 23772 274
rect 23716 220 23772 222
rect 23904 274 23960 276
rect 23904 222 23906 274
rect 23906 222 23958 274
rect 23958 222 23960 274
rect 23904 220 23960 222
rect 24964 274 25020 276
rect 24964 222 24966 274
rect 24966 222 25018 274
rect 25018 222 25020 274
rect 24964 220 25020 222
rect 25152 274 25208 276
rect 25152 222 25154 274
rect 25154 222 25206 274
rect 25206 222 25208 274
rect 25152 220 25208 222
rect 26212 274 26268 276
rect 26212 222 26214 274
rect 26214 222 26266 274
rect 26266 222 26268 274
rect 26212 220 26268 222
rect 26400 274 26456 276
rect 26400 222 26402 274
rect 26402 222 26454 274
rect 26454 222 26456 274
rect 26400 220 26456 222
rect 27460 274 27516 276
rect 27460 222 27462 274
rect 27462 222 27514 274
rect 27514 222 27516 274
rect 27460 220 27516 222
rect 27648 274 27704 276
rect 27648 222 27650 274
rect 27650 222 27702 274
rect 27702 222 27704 274
rect 27648 220 27704 222
rect 28708 274 28764 276
rect 28708 222 28710 274
rect 28710 222 28762 274
rect 28762 222 28764 274
rect 28708 220 28764 222
rect 28896 274 28952 276
rect 28896 222 28898 274
rect 28898 222 28950 274
rect 28950 222 28952 274
rect 28896 220 28952 222
rect 29956 274 30012 276
rect 29956 222 29958 274
rect 29958 222 30010 274
rect 30010 222 30012 274
rect 29956 220 30012 222
rect 30144 274 30200 276
rect 30144 222 30146 274
rect 30146 222 30198 274
rect 30198 222 30200 274
rect 30144 220 30200 222
rect 31204 274 31260 276
rect 31204 222 31206 274
rect 31206 222 31258 274
rect 31258 222 31260 274
rect 31204 220 31260 222
rect 31392 274 31448 276
rect 31392 222 31394 274
rect 31394 222 31446 274
rect 31446 222 31448 274
rect 31392 220 31448 222
rect 32452 274 32508 276
rect 32452 222 32454 274
rect 32454 222 32506 274
rect 32506 222 32508 274
rect 32452 220 32508 222
rect 32640 274 32696 276
rect 32640 222 32642 274
rect 32642 222 32694 274
rect 32694 222 32696 274
rect 32640 220 32696 222
rect 33700 274 33756 276
rect 33700 222 33702 274
rect 33702 222 33754 274
rect 33754 222 33756 274
rect 33700 220 33756 222
rect 33888 274 33944 276
rect 33888 222 33890 274
rect 33890 222 33942 274
rect 33942 222 33944 274
rect 33888 220 33944 222
rect 34948 274 35004 276
rect 34948 222 34950 274
rect 34950 222 35002 274
rect 35002 222 35004 274
rect 34948 220 35004 222
rect 35136 274 35192 276
rect 35136 222 35138 274
rect 35138 222 35190 274
rect 35190 222 35192 274
rect 35136 220 35192 222
rect 36196 274 36252 276
rect 36196 222 36198 274
rect 36198 222 36250 274
rect 36250 222 36252 274
rect 36196 220 36252 222
rect 36384 274 36440 276
rect 36384 222 36386 274
rect 36386 222 36438 274
rect 36438 222 36440 274
rect 36384 220 36440 222
rect 37444 274 37500 276
rect 37444 222 37446 274
rect 37446 222 37498 274
rect 37498 222 37500 274
rect 37444 220 37500 222
rect 37632 274 37688 276
rect 37632 222 37634 274
rect 37634 222 37686 274
rect 37686 222 37688 274
rect 37632 220 37688 222
rect 38692 274 38748 276
rect 38692 222 38694 274
rect 38694 222 38746 274
rect 38746 222 38748 274
rect 38692 220 38748 222
rect 38880 274 38936 276
rect 38880 222 38882 274
rect 38882 222 38934 274
rect 38934 222 38936 274
rect 38880 220 38936 222
rect 39940 274 39996 276
rect 39940 222 39942 274
rect 39942 222 39994 274
rect 39994 222 39996 274
rect 39940 220 39996 222
rect 40128 274 40184 276
rect 40128 222 40130 274
rect 40130 222 40182 274
rect 40182 222 40184 274
rect 40128 220 40184 222
rect 41188 274 41244 276
rect 41188 222 41190 274
rect 41190 222 41242 274
rect 41242 222 41244 274
rect 41188 220 41244 222
rect 41376 274 41432 276
rect 41376 222 41378 274
rect 41378 222 41430 274
rect 41430 222 41432 274
rect 41376 220 41432 222
rect 42436 274 42492 276
rect 42436 222 42438 274
rect 42438 222 42490 274
rect 42490 222 42492 274
rect 42436 220 42492 222
rect 42624 274 42680 276
rect 42624 222 42626 274
rect 42626 222 42678 274
rect 42678 222 42680 274
rect 42624 220 42680 222
rect 43684 274 43740 276
rect 43684 222 43686 274
rect 43686 222 43738 274
rect 43738 222 43740 274
rect 43684 220 43740 222
rect 43872 274 43928 276
rect 43872 222 43874 274
rect 43874 222 43926 274
rect 43926 222 43928 274
rect 43872 220 43928 222
rect 44932 274 44988 276
rect 44932 222 44934 274
rect 44934 222 44986 274
rect 44986 222 44988 274
rect 44932 220 44988 222
rect 45120 274 45176 276
rect 45120 222 45122 274
rect 45122 222 45174 274
rect 45174 222 45176 274
rect 45120 220 45176 222
rect 46180 274 46236 276
rect 46180 222 46182 274
rect 46182 222 46234 274
rect 46234 222 46236 274
rect 46180 220 46236 222
rect 46368 274 46424 276
rect 46368 222 46370 274
rect 46370 222 46422 274
rect 46422 222 46424 274
rect 46368 220 46424 222
rect 47428 274 47484 276
rect 47428 222 47430 274
rect 47430 222 47482 274
rect 47482 222 47484 274
rect 47428 220 47484 222
rect 47616 274 47672 276
rect 47616 222 47618 274
rect 47618 222 47670 274
rect 47670 222 47672 274
rect 47616 220 47672 222
rect 48676 274 48732 276
rect 48676 222 48678 274
rect 48678 222 48730 274
rect 48730 222 48732 274
rect 48676 220 48732 222
rect 48864 274 48920 276
rect 48864 222 48866 274
rect 48866 222 48918 274
rect 48918 222 48920 274
rect 48864 220 48920 222
rect 49924 274 49980 276
rect 49924 222 49926 274
rect 49926 222 49978 274
rect 49978 222 49980 274
rect 49924 220 49980 222
rect 50112 274 50168 276
rect 50112 222 50114 274
rect 50114 222 50166 274
rect 50166 222 50168 274
rect 50112 220 50168 222
rect 51172 274 51228 276
rect 51172 222 51174 274
rect 51174 222 51226 274
rect 51226 222 51228 274
rect 51172 220 51228 222
rect 51360 274 51416 276
rect 51360 222 51362 274
rect 51362 222 51414 274
rect 51414 222 51416 274
rect 51360 220 51416 222
rect 52420 274 52476 276
rect 52420 222 52422 274
rect 52422 222 52474 274
rect 52474 222 52476 274
rect 52420 220 52476 222
rect 52608 274 52664 276
rect 52608 222 52610 274
rect 52610 222 52662 274
rect 52662 222 52664 274
rect 52608 220 52664 222
rect 53668 274 53724 276
rect 53668 222 53670 274
rect 53670 222 53722 274
rect 53722 222 53724 274
rect 53668 220 53724 222
rect 53856 274 53912 276
rect 53856 222 53858 274
rect 53858 222 53910 274
rect 53910 222 53912 274
rect 53856 220 53912 222
rect 54916 274 54972 276
rect 54916 222 54918 274
rect 54918 222 54970 274
rect 54970 222 54972 274
rect 54916 220 54972 222
rect 55104 274 55160 276
rect 55104 222 55106 274
rect 55106 222 55158 274
rect 55158 222 55160 274
rect 55104 220 55160 222
rect 56164 274 56220 276
rect 56164 222 56166 274
rect 56166 222 56218 274
rect 56218 222 56220 274
rect 56164 220 56220 222
rect 56352 274 56408 276
rect 56352 222 56354 274
rect 56354 222 56406 274
rect 56406 222 56408 274
rect 56352 220 56408 222
rect 57412 274 57468 276
rect 57412 222 57414 274
rect 57414 222 57466 274
rect 57466 222 57468 274
rect 57412 220 57468 222
rect 57600 274 57656 276
rect 57600 222 57602 274
rect 57602 222 57654 274
rect 57654 222 57656 274
rect 57600 220 57656 222
rect 58660 274 58716 276
rect 58660 222 58662 274
rect 58662 222 58714 274
rect 58714 222 58716 274
rect 58660 220 58716 222
rect 58848 274 58904 276
rect 58848 222 58850 274
rect 58850 222 58902 274
rect 58902 222 58904 274
rect 58848 220 58904 222
rect 59908 274 59964 276
rect 59908 222 59910 274
rect 59910 222 59962 274
rect 59962 222 59964 274
rect 59908 220 59964 222
rect 60096 274 60152 276
rect 60096 222 60098 274
rect 60098 222 60150 274
rect 60150 222 60152 274
rect 60096 220 60152 222
rect 61156 274 61212 276
rect 61156 222 61158 274
rect 61158 222 61210 274
rect 61210 222 61212 274
rect 61156 220 61212 222
rect 61344 274 61400 276
rect 61344 222 61346 274
rect 61346 222 61398 274
rect 61398 222 61400 274
rect 61344 220 61400 222
rect 62404 274 62460 276
rect 62404 222 62406 274
rect 62406 222 62458 274
rect 62458 222 62460 274
rect 62404 220 62460 222
rect 62592 274 62648 276
rect 62592 222 62594 274
rect 62594 222 62646 274
rect 62646 222 62648 274
rect 62592 220 62648 222
rect 63652 274 63708 276
rect 63652 222 63654 274
rect 63654 222 63706 274
rect 63706 222 63708 274
rect 63652 220 63708 222
rect 63840 274 63896 276
rect 63840 222 63842 274
rect 63842 222 63894 274
rect 63894 222 63896 274
rect 63840 220 63896 222
rect 64900 274 64956 276
rect 64900 222 64902 274
rect 64902 222 64954 274
rect 64954 222 64956 274
rect 64900 220 64956 222
rect 65088 274 65144 276
rect 65088 222 65090 274
rect 65090 222 65142 274
rect 65142 222 65144 274
rect 65088 220 65144 222
rect 66148 274 66204 276
rect 66148 222 66150 274
rect 66150 222 66202 274
rect 66202 222 66204 274
rect 66148 220 66204 222
rect 66336 274 66392 276
rect 66336 222 66338 274
rect 66338 222 66390 274
rect 66390 222 66392 274
rect 66336 220 66392 222
rect 67396 274 67452 276
rect 67396 222 67398 274
rect 67398 222 67450 274
rect 67450 222 67452 274
rect 67396 220 67452 222
rect 67584 274 67640 276
rect 67584 222 67586 274
rect 67586 222 67638 274
rect 67638 222 67640 274
rect 67584 220 67640 222
rect 68644 274 68700 276
rect 68644 222 68646 274
rect 68646 222 68698 274
rect 68698 222 68700 274
rect 68644 220 68700 222
rect 68832 274 68888 276
rect 68832 222 68834 274
rect 68834 222 68886 274
rect 68886 222 68888 274
rect 68832 220 68888 222
rect 69892 274 69948 276
rect 69892 222 69894 274
rect 69894 222 69946 274
rect 69946 222 69948 274
rect 69892 220 69948 222
rect 70080 274 70136 276
rect 70080 222 70082 274
rect 70082 222 70134 274
rect 70134 222 70136 274
rect 70080 220 70136 222
rect 71140 274 71196 276
rect 71140 222 71142 274
rect 71142 222 71194 274
rect 71194 222 71196 274
rect 71140 220 71196 222
rect 71328 274 71384 276
rect 71328 222 71330 274
rect 71330 222 71382 274
rect 71382 222 71384 274
rect 71328 220 71384 222
rect 72388 274 72444 276
rect 72388 222 72390 274
rect 72390 222 72442 274
rect 72442 222 72444 274
rect 72388 220 72444 222
rect 72576 274 72632 276
rect 72576 222 72578 274
rect 72578 222 72630 274
rect 72630 222 72632 274
rect 72576 220 72632 222
rect 73636 274 73692 276
rect 73636 222 73638 274
rect 73638 222 73690 274
rect 73690 222 73692 274
rect 73636 220 73692 222
rect 73824 274 73880 276
rect 73824 222 73826 274
rect 73826 222 73878 274
rect 73878 222 73880 274
rect 73824 220 73880 222
rect 74884 274 74940 276
rect 74884 222 74886 274
rect 74886 222 74938 274
rect 74938 222 74940 274
rect 74884 220 74940 222
rect 75072 274 75128 276
rect 75072 222 75074 274
rect 75074 222 75126 274
rect 75126 222 75128 274
rect 75072 220 75128 222
rect 76132 274 76188 276
rect 76132 222 76134 274
rect 76134 222 76186 274
rect 76186 222 76188 274
rect 76132 220 76188 222
rect 76320 274 76376 276
rect 76320 222 76322 274
rect 76322 222 76374 274
rect 76374 222 76376 274
rect 76320 220 76376 222
rect 77380 274 77436 276
rect 77380 222 77382 274
rect 77382 222 77434 274
rect 77434 222 77436 274
rect 77380 220 77436 222
rect 77568 274 77624 276
rect 77568 222 77570 274
rect 77570 222 77622 274
rect 77622 222 77624 274
rect 77568 220 77624 222
rect 78628 274 78684 276
rect 78628 222 78630 274
rect 78630 222 78682 274
rect 78682 222 78684 274
rect 78628 220 78684 222
rect 78816 274 78872 276
rect 78816 222 78818 274
rect 78818 222 78870 274
rect 78870 222 78872 274
rect 78816 220 78872 222
rect 79876 274 79932 276
rect 79876 222 79878 274
rect 79878 222 79930 274
rect 79930 222 79932 274
rect 79876 220 79932 222
rect 80064 274 80120 276
rect 80064 222 80066 274
rect 80066 222 80118 274
rect 80118 222 80120 274
rect 80064 220 80120 222
rect 81124 274 81180 276
rect 81124 222 81126 274
rect 81126 222 81178 274
rect 81178 222 81180 274
rect 81124 220 81180 222
rect 1904 150 1960 152
rect 1904 98 1906 150
rect 1906 98 1958 150
rect 1958 98 1960 150
rect 1904 96 1960 98
rect 2036 150 2092 152
rect 2036 98 2038 150
rect 2038 98 2090 150
rect 2090 98 2092 150
rect 2036 96 2092 98
rect 3152 150 3208 152
rect 3152 98 3154 150
rect 3154 98 3206 150
rect 3206 98 3208 150
rect 3152 96 3208 98
rect 3284 150 3340 152
rect 3284 98 3286 150
rect 3286 98 3338 150
rect 3338 98 3340 150
rect 3284 96 3340 98
rect 4400 150 4456 152
rect 4400 98 4402 150
rect 4402 98 4454 150
rect 4454 98 4456 150
rect 4400 96 4456 98
rect 4532 150 4588 152
rect 4532 98 4534 150
rect 4534 98 4586 150
rect 4586 98 4588 150
rect 4532 96 4588 98
rect 5648 150 5704 152
rect 5648 98 5650 150
rect 5650 98 5702 150
rect 5702 98 5704 150
rect 5648 96 5704 98
rect 5780 150 5836 152
rect 5780 98 5782 150
rect 5782 98 5834 150
rect 5834 98 5836 150
rect 5780 96 5836 98
rect 6896 150 6952 152
rect 6896 98 6898 150
rect 6898 98 6950 150
rect 6950 98 6952 150
rect 6896 96 6952 98
rect 7028 150 7084 152
rect 7028 98 7030 150
rect 7030 98 7082 150
rect 7082 98 7084 150
rect 7028 96 7084 98
rect 8144 150 8200 152
rect 8144 98 8146 150
rect 8146 98 8198 150
rect 8198 98 8200 150
rect 8144 96 8200 98
rect 8276 150 8332 152
rect 8276 98 8278 150
rect 8278 98 8330 150
rect 8330 98 8332 150
rect 8276 96 8332 98
rect 9392 150 9448 152
rect 9392 98 9394 150
rect 9394 98 9446 150
rect 9446 98 9448 150
rect 9392 96 9448 98
rect 9524 150 9580 152
rect 9524 98 9526 150
rect 9526 98 9578 150
rect 9578 98 9580 150
rect 9524 96 9580 98
rect 10640 150 10696 152
rect 10640 98 10642 150
rect 10642 98 10694 150
rect 10694 98 10696 150
rect 10640 96 10696 98
rect 10772 150 10828 152
rect 10772 98 10774 150
rect 10774 98 10826 150
rect 10826 98 10828 150
rect 10772 96 10828 98
rect 11888 150 11944 152
rect 11888 98 11890 150
rect 11890 98 11942 150
rect 11942 98 11944 150
rect 11888 96 11944 98
rect 12020 150 12076 152
rect 12020 98 12022 150
rect 12022 98 12074 150
rect 12074 98 12076 150
rect 12020 96 12076 98
rect 13136 150 13192 152
rect 13136 98 13138 150
rect 13138 98 13190 150
rect 13190 98 13192 150
rect 13136 96 13192 98
rect 13268 150 13324 152
rect 13268 98 13270 150
rect 13270 98 13322 150
rect 13322 98 13324 150
rect 13268 96 13324 98
rect 14384 150 14440 152
rect 14384 98 14386 150
rect 14386 98 14438 150
rect 14438 98 14440 150
rect 14384 96 14440 98
rect 14516 150 14572 152
rect 14516 98 14518 150
rect 14518 98 14570 150
rect 14570 98 14572 150
rect 14516 96 14572 98
rect 15632 150 15688 152
rect 15632 98 15634 150
rect 15634 98 15686 150
rect 15686 98 15688 150
rect 15632 96 15688 98
rect 15764 150 15820 152
rect 15764 98 15766 150
rect 15766 98 15818 150
rect 15818 98 15820 150
rect 15764 96 15820 98
rect 16880 150 16936 152
rect 16880 98 16882 150
rect 16882 98 16934 150
rect 16934 98 16936 150
rect 16880 96 16936 98
rect 17012 150 17068 152
rect 17012 98 17014 150
rect 17014 98 17066 150
rect 17066 98 17068 150
rect 17012 96 17068 98
rect 18128 150 18184 152
rect 18128 98 18130 150
rect 18130 98 18182 150
rect 18182 98 18184 150
rect 18128 96 18184 98
rect 18260 150 18316 152
rect 18260 98 18262 150
rect 18262 98 18314 150
rect 18314 98 18316 150
rect 18260 96 18316 98
rect 19376 150 19432 152
rect 19376 98 19378 150
rect 19378 98 19430 150
rect 19430 98 19432 150
rect 19376 96 19432 98
rect 19508 150 19564 152
rect 19508 98 19510 150
rect 19510 98 19562 150
rect 19562 98 19564 150
rect 19508 96 19564 98
rect 20624 150 20680 152
rect 20624 98 20626 150
rect 20626 98 20678 150
rect 20678 98 20680 150
rect 20624 96 20680 98
rect 20756 150 20812 152
rect 20756 98 20758 150
rect 20758 98 20810 150
rect 20810 98 20812 150
rect 20756 96 20812 98
rect 21872 150 21928 152
rect 21872 98 21874 150
rect 21874 98 21926 150
rect 21926 98 21928 150
rect 21872 96 21928 98
rect 22004 150 22060 152
rect 22004 98 22006 150
rect 22006 98 22058 150
rect 22058 98 22060 150
rect 22004 96 22060 98
rect 23120 150 23176 152
rect 23120 98 23122 150
rect 23122 98 23174 150
rect 23174 98 23176 150
rect 23120 96 23176 98
rect 23252 150 23308 152
rect 23252 98 23254 150
rect 23254 98 23306 150
rect 23306 98 23308 150
rect 23252 96 23308 98
rect 24368 150 24424 152
rect 24368 98 24370 150
rect 24370 98 24422 150
rect 24422 98 24424 150
rect 24368 96 24424 98
rect 24500 150 24556 152
rect 24500 98 24502 150
rect 24502 98 24554 150
rect 24554 98 24556 150
rect 24500 96 24556 98
rect 25616 150 25672 152
rect 25616 98 25618 150
rect 25618 98 25670 150
rect 25670 98 25672 150
rect 25616 96 25672 98
rect 25748 150 25804 152
rect 25748 98 25750 150
rect 25750 98 25802 150
rect 25802 98 25804 150
rect 25748 96 25804 98
rect 26864 150 26920 152
rect 26864 98 26866 150
rect 26866 98 26918 150
rect 26918 98 26920 150
rect 26864 96 26920 98
rect 26996 150 27052 152
rect 26996 98 26998 150
rect 26998 98 27050 150
rect 27050 98 27052 150
rect 26996 96 27052 98
rect 28112 150 28168 152
rect 28112 98 28114 150
rect 28114 98 28166 150
rect 28166 98 28168 150
rect 28112 96 28168 98
rect 28244 150 28300 152
rect 28244 98 28246 150
rect 28246 98 28298 150
rect 28298 98 28300 150
rect 28244 96 28300 98
rect 29360 150 29416 152
rect 29360 98 29362 150
rect 29362 98 29414 150
rect 29414 98 29416 150
rect 29360 96 29416 98
rect 29492 150 29548 152
rect 29492 98 29494 150
rect 29494 98 29546 150
rect 29546 98 29548 150
rect 29492 96 29548 98
rect 30608 150 30664 152
rect 30608 98 30610 150
rect 30610 98 30662 150
rect 30662 98 30664 150
rect 30608 96 30664 98
rect 30740 150 30796 152
rect 30740 98 30742 150
rect 30742 98 30794 150
rect 30794 98 30796 150
rect 30740 96 30796 98
rect 31856 150 31912 152
rect 31856 98 31858 150
rect 31858 98 31910 150
rect 31910 98 31912 150
rect 31856 96 31912 98
rect 31988 150 32044 152
rect 31988 98 31990 150
rect 31990 98 32042 150
rect 32042 98 32044 150
rect 31988 96 32044 98
rect 33104 150 33160 152
rect 33104 98 33106 150
rect 33106 98 33158 150
rect 33158 98 33160 150
rect 33104 96 33160 98
rect 33236 150 33292 152
rect 33236 98 33238 150
rect 33238 98 33290 150
rect 33290 98 33292 150
rect 33236 96 33292 98
rect 34352 150 34408 152
rect 34352 98 34354 150
rect 34354 98 34406 150
rect 34406 98 34408 150
rect 34352 96 34408 98
rect 34484 150 34540 152
rect 34484 98 34486 150
rect 34486 98 34538 150
rect 34538 98 34540 150
rect 34484 96 34540 98
rect 35600 150 35656 152
rect 35600 98 35602 150
rect 35602 98 35654 150
rect 35654 98 35656 150
rect 35600 96 35656 98
rect 35732 150 35788 152
rect 35732 98 35734 150
rect 35734 98 35786 150
rect 35786 98 35788 150
rect 35732 96 35788 98
rect 36848 150 36904 152
rect 36848 98 36850 150
rect 36850 98 36902 150
rect 36902 98 36904 150
rect 36848 96 36904 98
rect 36980 150 37036 152
rect 36980 98 36982 150
rect 36982 98 37034 150
rect 37034 98 37036 150
rect 36980 96 37036 98
rect 38096 150 38152 152
rect 38096 98 38098 150
rect 38098 98 38150 150
rect 38150 98 38152 150
rect 38096 96 38152 98
rect 38228 150 38284 152
rect 38228 98 38230 150
rect 38230 98 38282 150
rect 38282 98 38284 150
rect 38228 96 38284 98
rect 39344 150 39400 152
rect 39344 98 39346 150
rect 39346 98 39398 150
rect 39398 98 39400 150
rect 39344 96 39400 98
rect 39476 150 39532 152
rect 39476 98 39478 150
rect 39478 98 39530 150
rect 39530 98 39532 150
rect 39476 96 39532 98
rect 40592 150 40648 152
rect 40592 98 40594 150
rect 40594 98 40646 150
rect 40646 98 40648 150
rect 40592 96 40648 98
rect 40724 150 40780 152
rect 40724 98 40726 150
rect 40726 98 40778 150
rect 40778 98 40780 150
rect 40724 96 40780 98
rect 41840 150 41896 152
rect 41840 98 41842 150
rect 41842 98 41894 150
rect 41894 98 41896 150
rect 41840 96 41896 98
rect 41972 150 42028 152
rect 41972 98 41974 150
rect 41974 98 42026 150
rect 42026 98 42028 150
rect 41972 96 42028 98
rect 43088 150 43144 152
rect 43088 98 43090 150
rect 43090 98 43142 150
rect 43142 98 43144 150
rect 43088 96 43144 98
rect 43220 150 43276 152
rect 43220 98 43222 150
rect 43222 98 43274 150
rect 43274 98 43276 150
rect 43220 96 43276 98
rect 44336 150 44392 152
rect 44336 98 44338 150
rect 44338 98 44390 150
rect 44390 98 44392 150
rect 44336 96 44392 98
rect 44468 150 44524 152
rect 44468 98 44470 150
rect 44470 98 44522 150
rect 44522 98 44524 150
rect 44468 96 44524 98
rect 45584 150 45640 152
rect 45584 98 45586 150
rect 45586 98 45638 150
rect 45638 98 45640 150
rect 45584 96 45640 98
rect 45716 150 45772 152
rect 45716 98 45718 150
rect 45718 98 45770 150
rect 45770 98 45772 150
rect 45716 96 45772 98
rect 46832 150 46888 152
rect 46832 98 46834 150
rect 46834 98 46886 150
rect 46886 98 46888 150
rect 46832 96 46888 98
rect 46964 150 47020 152
rect 46964 98 46966 150
rect 46966 98 47018 150
rect 47018 98 47020 150
rect 46964 96 47020 98
rect 48080 150 48136 152
rect 48080 98 48082 150
rect 48082 98 48134 150
rect 48134 98 48136 150
rect 48080 96 48136 98
rect 48212 150 48268 152
rect 48212 98 48214 150
rect 48214 98 48266 150
rect 48266 98 48268 150
rect 48212 96 48268 98
rect 49328 150 49384 152
rect 49328 98 49330 150
rect 49330 98 49382 150
rect 49382 98 49384 150
rect 49328 96 49384 98
rect 49460 150 49516 152
rect 49460 98 49462 150
rect 49462 98 49514 150
rect 49514 98 49516 150
rect 49460 96 49516 98
rect 50576 150 50632 152
rect 50576 98 50578 150
rect 50578 98 50630 150
rect 50630 98 50632 150
rect 50576 96 50632 98
rect 50708 150 50764 152
rect 50708 98 50710 150
rect 50710 98 50762 150
rect 50762 98 50764 150
rect 50708 96 50764 98
rect 51824 150 51880 152
rect 51824 98 51826 150
rect 51826 98 51878 150
rect 51878 98 51880 150
rect 51824 96 51880 98
rect 51956 150 52012 152
rect 51956 98 51958 150
rect 51958 98 52010 150
rect 52010 98 52012 150
rect 51956 96 52012 98
rect 53072 150 53128 152
rect 53072 98 53074 150
rect 53074 98 53126 150
rect 53126 98 53128 150
rect 53072 96 53128 98
rect 53204 150 53260 152
rect 53204 98 53206 150
rect 53206 98 53258 150
rect 53258 98 53260 150
rect 53204 96 53260 98
rect 54320 150 54376 152
rect 54320 98 54322 150
rect 54322 98 54374 150
rect 54374 98 54376 150
rect 54320 96 54376 98
rect 54452 150 54508 152
rect 54452 98 54454 150
rect 54454 98 54506 150
rect 54506 98 54508 150
rect 54452 96 54508 98
rect 55568 150 55624 152
rect 55568 98 55570 150
rect 55570 98 55622 150
rect 55622 98 55624 150
rect 55568 96 55624 98
rect 55700 150 55756 152
rect 55700 98 55702 150
rect 55702 98 55754 150
rect 55754 98 55756 150
rect 55700 96 55756 98
rect 56816 150 56872 152
rect 56816 98 56818 150
rect 56818 98 56870 150
rect 56870 98 56872 150
rect 56816 96 56872 98
rect 56948 150 57004 152
rect 56948 98 56950 150
rect 56950 98 57002 150
rect 57002 98 57004 150
rect 56948 96 57004 98
rect 58064 150 58120 152
rect 58064 98 58066 150
rect 58066 98 58118 150
rect 58118 98 58120 150
rect 58064 96 58120 98
rect 58196 150 58252 152
rect 58196 98 58198 150
rect 58198 98 58250 150
rect 58250 98 58252 150
rect 58196 96 58252 98
rect 59312 150 59368 152
rect 59312 98 59314 150
rect 59314 98 59366 150
rect 59366 98 59368 150
rect 59312 96 59368 98
rect 59444 150 59500 152
rect 59444 98 59446 150
rect 59446 98 59498 150
rect 59498 98 59500 150
rect 59444 96 59500 98
rect 60560 150 60616 152
rect 60560 98 60562 150
rect 60562 98 60614 150
rect 60614 98 60616 150
rect 60560 96 60616 98
rect 60692 150 60748 152
rect 60692 98 60694 150
rect 60694 98 60746 150
rect 60746 98 60748 150
rect 60692 96 60748 98
rect 61808 150 61864 152
rect 61808 98 61810 150
rect 61810 98 61862 150
rect 61862 98 61864 150
rect 61808 96 61864 98
rect 61940 150 61996 152
rect 61940 98 61942 150
rect 61942 98 61994 150
rect 61994 98 61996 150
rect 61940 96 61996 98
rect 63056 150 63112 152
rect 63056 98 63058 150
rect 63058 98 63110 150
rect 63110 98 63112 150
rect 63056 96 63112 98
rect 63188 150 63244 152
rect 63188 98 63190 150
rect 63190 98 63242 150
rect 63242 98 63244 150
rect 63188 96 63244 98
rect 64304 150 64360 152
rect 64304 98 64306 150
rect 64306 98 64358 150
rect 64358 98 64360 150
rect 64304 96 64360 98
rect 64436 150 64492 152
rect 64436 98 64438 150
rect 64438 98 64490 150
rect 64490 98 64492 150
rect 64436 96 64492 98
rect 65552 150 65608 152
rect 65552 98 65554 150
rect 65554 98 65606 150
rect 65606 98 65608 150
rect 65552 96 65608 98
rect 65684 150 65740 152
rect 65684 98 65686 150
rect 65686 98 65738 150
rect 65738 98 65740 150
rect 65684 96 65740 98
rect 66800 150 66856 152
rect 66800 98 66802 150
rect 66802 98 66854 150
rect 66854 98 66856 150
rect 66800 96 66856 98
rect 66932 150 66988 152
rect 66932 98 66934 150
rect 66934 98 66986 150
rect 66986 98 66988 150
rect 66932 96 66988 98
rect 68048 150 68104 152
rect 68048 98 68050 150
rect 68050 98 68102 150
rect 68102 98 68104 150
rect 68048 96 68104 98
rect 68180 150 68236 152
rect 68180 98 68182 150
rect 68182 98 68234 150
rect 68234 98 68236 150
rect 68180 96 68236 98
rect 69296 150 69352 152
rect 69296 98 69298 150
rect 69298 98 69350 150
rect 69350 98 69352 150
rect 69296 96 69352 98
rect 69428 150 69484 152
rect 69428 98 69430 150
rect 69430 98 69482 150
rect 69482 98 69484 150
rect 69428 96 69484 98
rect 70544 150 70600 152
rect 70544 98 70546 150
rect 70546 98 70598 150
rect 70598 98 70600 150
rect 70544 96 70600 98
rect 70676 150 70732 152
rect 70676 98 70678 150
rect 70678 98 70730 150
rect 70730 98 70732 150
rect 70676 96 70732 98
rect 71792 150 71848 152
rect 71792 98 71794 150
rect 71794 98 71846 150
rect 71846 98 71848 150
rect 71792 96 71848 98
rect 71924 150 71980 152
rect 71924 98 71926 150
rect 71926 98 71978 150
rect 71978 98 71980 150
rect 71924 96 71980 98
rect 73040 150 73096 152
rect 73040 98 73042 150
rect 73042 98 73094 150
rect 73094 98 73096 150
rect 73040 96 73096 98
rect 73172 150 73228 152
rect 73172 98 73174 150
rect 73174 98 73226 150
rect 73226 98 73228 150
rect 73172 96 73228 98
rect 74288 150 74344 152
rect 74288 98 74290 150
rect 74290 98 74342 150
rect 74342 98 74344 150
rect 74288 96 74344 98
rect 74420 150 74476 152
rect 74420 98 74422 150
rect 74422 98 74474 150
rect 74474 98 74476 150
rect 74420 96 74476 98
rect 75536 150 75592 152
rect 75536 98 75538 150
rect 75538 98 75590 150
rect 75590 98 75592 150
rect 75536 96 75592 98
rect 75668 150 75724 152
rect 75668 98 75670 150
rect 75670 98 75722 150
rect 75722 98 75724 150
rect 75668 96 75724 98
rect 76784 150 76840 152
rect 76784 98 76786 150
rect 76786 98 76838 150
rect 76838 98 76840 150
rect 76784 96 76840 98
rect 76916 150 76972 152
rect 76916 98 76918 150
rect 76918 98 76970 150
rect 76970 98 76972 150
rect 76916 96 76972 98
rect 78032 150 78088 152
rect 78032 98 78034 150
rect 78034 98 78086 150
rect 78086 98 78088 150
rect 78032 96 78088 98
rect 78164 150 78220 152
rect 78164 98 78166 150
rect 78166 98 78218 150
rect 78218 98 78220 150
rect 78164 96 78220 98
rect 79280 150 79336 152
rect 79280 98 79282 150
rect 79282 98 79334 150
rect 79334 98 79336 150
rect 79280 96 79336 98
rect 79412 150 79468 152
rect 79412 98 79414 150
rect 79414 98 79466 150
rect 79466 98 79468 150
rect 79412 96 79468 98
rect 80528 150 80584 152
rect 80528 98 80530 150
rect 80530 98 80582 150
rect 80582 98 80584 150
rect 80528 96 80584 98
rect 80660 150 80716 152
rect 80660 98 80662 150
rect 80662 98 80714 150
rect 80714 98 80716 150
rect 80660 96 80716 98
<< metal3 >>
rect 1949 1482 2047 1580
rect 3197 1482 3295 1580
rect 4445 1482 4543 1580
rect 5693 1482 5791 1580
rect 6941 1482 7039 1580
rect 8189 1482 8287 1580
rect 9437 1482 9535 1580
rect 10685 1482 10783 1580
rect 11933 1482 12031 1580
rect 13181 1482 13279 1580
rect 14429 1482 14527 1580
rect 15677 1482 15775 1580
rect 16925 1482 17023 1580
rect 18173 1482 18271 1580
rect 19421 1482 19519 1580
rect 20669 1482 20767 1580
rect 21917 1482 22015 1580
rect 23165 1482 23263 1580
rect 24413 1482 24511 1580
rect 25661 1482 25759 1580
rect 26909 1482 27007 1580
rect 28157 1482 28255 1580
rect 29405 1482 29503 1580
rect 30653 1482 30751 1580
rect 31901 1482 31999 1580
rect 33149 1482 33247 1580
rect 34397 1482 34495 1580
rect 35645 1482 35743 1580
rect 36893 1482 36991 1580
rect 38141 1482 38239 1580
rect 39389 1482 39487 1580
rect 40637 1482 40735 1580
rect 41885 1482 41983 1580
rect 43133 1482 43231 1580
rect 44381 1482 44479 1580
rect 45629 1482 45727 1580
rect 46877 1482 46975 1580
rect 48125 1482 48223 1580
rect 49373 1482 49471 1580
rect 50621 1482 50719 1580
rect 51869 1482 51967 1580
rect 53117 1482 53215 1580
rect 54365 1482 54463 1580
rect 55613 1482 55711 1580
rect 56861 1482 56959 1580
rect 58109 1482 58207 1580
rect 59357 1482 59455 1580
rect 60605 1482 60703 1580
rect 61853 1482 61951 1580
rect 63101 1482 63199 1580
rect 64349 1482 64447 1580
rect 65597 1482 65695 1580
rect 66845 1482 66943 1580
rect 68093 1482 68191 1580
rect 69341 1482 69439 1580
rect 70589 1482 70687 1580
rect 71837 1482 71935 1580
rect 73085 1482 73183 1580
rect 74333 1482 74431 1580
rect 75581 1482 75679 1580
rect 76829 1482 76927 1580
rect 78077 1482 78175 1580
rect 79325 1482 79423 1580
rect 80573 1482 80671 1580
rect 3525 804 3591 807
rect 6021 804 6087 807
rect 8517 804 8583 807
rect 11013 804 11079 807
rect 13509 804 13575 807
rect 16005 804 16071 807
rect 18501 804 18567 807
rect 20997 804 21063 807
rect 23493 804 23559 807
rect 25989 804 26055 807
rect 28485 804 28551 807
rect 30981 804 31047 807
rect 33477 804 33543 807
rect 35973 804 36039 807
rect 38469 804 38535 807
rect 40965 804 41031 807
rect 43461 804 43527 807
rect 45957 804 46023 807
rect 48453 804 48519 807
rect 50949 804 51015 807
rect 53445 804 53511 807
rect 55941 804 56007 807
rect 58437 804 58503 807
rect 60933 804 60999 807
rect 63429 804 63495 807
rect 65925 804 65991 807
rect 68421 804 68487 807
rect 70917 804 70983 807
rect 73413 804 73479 807
rect 75909 804 75975 807
rect 78405 804 78471 807
rect 80901 804 80967 807
rect 0 802 81246 804
rect 0 746 3530 802
rect 3586 746 6026 802
rect 6082 746 8522 802
rect 8578 746 11018 802
rect 11074 746 13514 802
rect 13570 746 16010 802
rect 16066 746 18506 802
rect 18562 746 21002 802
rect 21058 746 23498 802
rect 23554 746 25994 802
rect 26050 746 28490 802
rect 28546 746 30986 802
rect 31042 746 33482 802
rect 33538 746 35978 802
rect 36034 746 38474 802
rect 38530 746 40970 802
rect 41026 746 43466 802
rect 43522 746 45962 802
rect 46018 746 48458 802
rect 48514 746 50954 802
rect 51010 746 53450 802
rect 53506 746 55946 802
rect 56002 746 58442 802
rect 58498 746 60938 802
rect 60994 746 63434 802
rect 63490 746 65930 802
rect 65986 746 68426 802
rect 68482 746 70922 802
rect 70978 746 73418 802
rect 73474 746 75914 802
rect 75970 746 78410 802
rect 78466 746 80906 802
rect 80962 746 81246 802
rect 0 744 81246 746
rect 3525 741 3591 744
rect 6021 741 6087 744
rect 8517 741 8583 744
rect 11013 741 11079 744
rect 13509 741 13575 744
rect 16005 741 16071 744
rect 18501 741 18567 744
rect 20997 741 21063 744
rect 23493 741 23559 744
rect 25989 741 26055 744
rect 28485 741 28551 744
rect 30981 741 31047 744
rect 33477 741 33543 744
rect 35973 741 36039 744
rect 38469 741 38535 744
rect 40965 741 41031 744
rect 43461 741 43527 744
rect 45957 741 46023 744
rect 48453 741 48519 744
rect 50949 741 51015 744
rect 53445 741 53511 744
rect 55941 741 56007 744
rect 58437 741 58503 744
rect 60933 741 60999 744
rect 63429 741 63495 744
rect 65925 741 65991 744
rect 68421 741 68487 744
rect 70917 741 70983 744
rect 73413 741 73479 744
rect 75909 741 75975 744
rect 78405 741 78471 744
rect 80901 741 80967 744
rect 2901 680 2967 683
rect 5397 680 5463 683
rect 7893 680 7959 683
rect 10389 680 10455 683
rect 12885 680 12951 683
rect 15381 680 15447 683
rect 17877 680 17943 683
rect 20373 680 20439 683
rect 22869 680 22935 683
rect 25365 680 25431 683
rect 27861 680 27927 683
rect 30357 680 30423 683
rect 32853 680 32919 683
rect 35349 680 35415 683
rect 37845 680 37911 683
rect 40341 680 40407 683
rect 42837 680 42903 683
rect 45333 680 45399 683
rect 47829 680 47895 683
rect 50325 680 50391 683
rect 52821 680 52887 683
rect 55317 680 55383 683
rect 57813 680 57879 683
rect 60309 680 60375 683
rect 62805 680 62871 683
rect 65301 680 65367 683
rect 67797 680 67863 683
rect 70293 680 70359 683
rect 72789 680 72855 683
rect 75285 680 75351 683
rect 77781 680 77847 683
rect 80277 680 80343 683
rect 0 678 81246 680
rect 0 622 2906 678
rect 2962 622 5402 678
rect 5458 622 7898 678
rect 7954 622 10394 678
rect 10450 622 12890 678
rect 12946 622 15386 678
rect 15442 622 17882 678
rect 17938 622 20378 678
rect 20434 622 22874 678
rect 22930 622 25370 678
rect 25426 622 27866 678
rect 27922 622 30362 678
rect 30418 622 32858 678
rect 32914 622 35354 678
rect 35410 622 37850 678
rect 37906 622 40346 678
rect 40402 622 42842 678
rect 42898 622 45338 678
rect 45394 622 47834 678
rect 47890 622 50330 678
rect 50386 622 52826 678
rect 52882 622 55322 678
rect 55378 622 57818 678
rect 57874 622 60314 678
rect 60370 622 62810 678
rect 62866 622 65306 678
rect 65362 622 67802 678
rect 67858 622 70298 678
rect 70354 622 72794 678
rect 72850 622 75290 678
rect 75346 622 77786 678
rect 77842 622 80282 678
rect 80338 622 81246 678
rect 0 620 81246 622
rect 2901 617 2967 620
rect 5397 617 5463 620
rect 7893 617 7959 620
rect 10389 617 10455 620
rect 12885 617 12951 620
rect 15381 617 15447 620
rect 17877 617 17943 620
rect 20373 617 20439 620
rect 22869 617 22935 620
rect 25365 617 25431 620
rect 27861 617 27927 620
rect 30357 617 30423 620
rect 32853 617 32919 620
rect 35349 617 35415 620
rect 37845 617 37911 620
rect 40341 617 40407 620
rect 42837 617 42903 620
rect 45333 617 45399 620
rect 47829 617 47895 620
rect 50325 617 50391 620
rect 52821 617 52887 620
rect 55317 617 55383 620
rect 57813 617 57879 620
rect 60309 617 60375 620
rect 62805 617 62871 620
rect 65301 617 65367 620
rect 67797 617 67863 620
rect 70293 617 70359 620
rect 72789 617 72855 620
rect 75285 617 75351 620
rect 77781 617 77847 620
rect 80277 617 80343 620
rect 2277 556 2343 559
rect 4773 556 4839 559
rect 7269 556 7335 559
rect 9765 556 9831 559
rect 12261 556 12327 559
rect 14757 556 14823 559
rect 17253 556 17319 559
rect 19749 556 19815 559
rect 22245 556 22311 559
rect 24741 556 24807 559
rect 27237 556 27303 559
rect 29733 556 29799 559
rect 32229 556 32295 559
rect 34725 556 34791 559
rect 37221 556 37287 559
rect 39717 556 39783 559
rect 42213 556 42279 559
rect 44709 556 44775 559
rect 47205 556 47271 559
rect 49701 556 49767 559
rect 52197 556 52263 559
rect 54693 556 54759 559
rect 57189 556 57255 559
rect 59685 556 59751 559
rect 62181 556 62247 559
rect 64677 556 64743 559
rect 67173 556 67239 559
rect 69669 556 69735 559
rect 72165 556 72231 559
rect 74661 556 74727 559
rect 77157 556 77223 559
rect 79653 556 79719 559
rect 0 554 81246 556
rect 0 498 2282 554
rect 2338 498 4778 554
rect 4834 498 7274 554
rect 7330 498 9770 554
rect 9826 498 12266 554
rect 12322 498 14762 554
rect 14818 498 17258 554
rect 17314 498 19754 554
rect 19810 498 22250 554
rect 22306 498 24746 554
rect 24802 498 27242 554
rect 27298 498 29738 554
rect 29794 498 32234 554
rect 32290 498 34730 554
rect 34786 498 37226 554
rect 37282 498 39722 554
rect 39778 498 42218 554
rect 42274 498 44714 554
rect 44770 498 47210 554
rect 47266 498 49706 554
rect 49762 498 52202 554
rect 52258 498 54698 554
rect 54754 498 57194 554
rect 57250 498 59690 554
rect 59746 498 62186 554
rect 62242 498 64682 554
rect 64738 498 67178 554
rect 67234 498 69674 554
rect 69730 498 72170 554
rect 72226 498 74666 554
rect 74722 498 77162 554
rect 77218 498 79658 554
rect 79714 498 81246 554
rect 0 496 81246 498
rect 2277 493 2343 496
rect 4773 493 4839 496
rect 7269 493 7335 496
rect 9765 493 9831 496
rect 12261 493 12327 496
rect 14757 493 14823 496
rect 17253 493 17319 496
rect 19749 493 19815 496
rect 22245 493 22311 496
rect 24741 493 24807 496
rect 27237 493 27303 496
rect 29733 493 29799 496
rect 32229 493 32295 496
rect 34725 493 34791 496
rect 37221 493 37287 496
rect 39717 493 39783 496
rect 42213 493 42279 496
rect 44709 493 44775 496
rect 47205 493 47271 496
rect 49701 493 49767 496
rect 52197 493 52263 496
rect 54693 493 54759 496
rect 57189 493 57255 496
rect 59685 493 59751 496
rect 62181 493 62247 496
rect 64677 493 64743 496
rect 67173 493 67239 496
rect 69669 493 69735 496
rect 72165 493 72231 496
rect 74661 493 74727 496
rect 77157 493 77223 496
rect 79653 493 79719 496
rect 1653 432 1719 435
rect 4149 432 4215 435
rect 6645 432 6711 435
rect 9141 432 9207 435
rect 11637 432 11703 435
rect 14133 432 14199 435
rect 16629 432 16695 435
rect 19125 432 19191 435
rect 21621 432 21687 435
rect 24117 432 24183 435
rect 26613 432 26679 435
rect 29109 432 29175 435
rect 31605 432 31671 435
rect 34101 432 34167 435
rect 36597 432 36663 435
rect 39093 432 39159 435
rect 41589 432 41655 435
rect 44085 432 44151 435
rect 46581 432 46647 435
rect 49077 432 49143 435
rect 51573 432 51639 435
rect 54069 432 54135 435
rect 56565 432 56631 435
rect 59061 432 59127 435
rect 61557 432 61623 435
rect 64053 432 64119 435
rect 66549 432 66615 435
rect 69045 432 69111 435
rect 71541 432 71607 435
rect 74037 432 74103 435
rect 76533 432 76599 435
rect 79029 432 79095 435
rect 0 430 81246 432
rect 0 374 1658 430
rect 1714 374 4154 430
rect 4210 374 6650 430
rect 6706 374 9146 430
rect 9202 374 11642 430
rect 11698 374 14138 430
rect 14194 374 16634 430
rect 16690 374 19130 430
rect 19186 374 21626 430
rect 21682 374 24122 430
rect 24178 374 26618 430
rect 26674 374 29114 430
rect 29170 374 31610 430
rect 31666 374 34106 430
rect 34162 374 36602 430
rect 36658 374 39098 430
rect 39154 374 41594 430
rect 41650 374 44090 430
rect 44146 374 46586 430
rect 46642 374 49082 430
rect 49138 374 51578 430
rect 51634 374 54074 430
rect 54130 374 56570 430
rect 56626 374 59066 430
rect 59122 374 61562 430
rect 61618 374 64058 430
rect 64114 374 66554 430
rect 66610 374 69050 430
rect 69106 374 71546 430
rect 71602 374 74042 430
rect 74098 374 76538 430
rect 76594 374 79034 430
rect 79090 374 81246 430
rect 0 372 81246 374
rect 1653 369 1719 372
rect 4149 369 4215 372
rect 6645 369 6711 372
rect 9141 369 9207 372
rect 11637 369 11703 372
rect 14133 369 14199 372
rect 16629 369 16695 372
rect 19125 369 19191 372
rect 21621 369 21687 372
rect 24117 369 24183 372
rect 26613 369 26679 372
rect 29109 369 29175 372
rect 31605 369 31671 372
rect 34101 369 34167 372
rect 36597 369 36663 372
rect 39093 369 39159 372
rect 41589 369 41655 372
rect 44085 369 44151 372
rect 46581 369 46647 372
rect 49077 369 49143 372
rect 51573 369 51639 372
rect 54069 369 54135 372
rect 56565 369 56631 372
rect 59061 369 59127 372
rect 61557 369 61623 372
rect 64053 369 64119 372
rect 66549 369 66615 372
rect 69045 369 69111 372
rect 71541 369 71607 372
rect 74037 369 74103 372
rect 76533 369 76599 372
rect 79029 369 79095 372
rect 1435 278 1501 281
rect 2495 278 2561 281
rect 2683 278 2749 281
rect 3743 278 3809 281
rect 1435 276 3809 278
rect 1435 220 1440 276
rect 1496 220 2500 276
rect 2556 220 2688 276
rect 2744 220 3748 276
rect 3804 220 3809 276
rect 1435 218 3809 220
rect 1435 215 1501 218
rect 2495 215 2561 218
rect 2683 215 2749 218
rect 3743 215 3809 218
rect 3931 278 3997 281
rect 4991 278 5057 281
rect 5179 278 5245 281
rect 6239 278 6305 281
rect 3931 276 6305 278
rect 3931 220 3936 276
rect 3992 220 4996 276
rect 5052 220 5184 276
rect 5240 220 6244 276
rect 6300 220 6305 276
rect 3931 218 6305 220
rect 3931 215 3997 218
rect 4991 215 5057 218
rect 5179 215 5245 218
rect 6239 215 6305 218
rect 6427 278 6493 281
rect 7487 278 7553 281
rect 7675 278 7741 281
rect 8735 278 8801 281
rect 6427 276 8801 278
rect 6427 220 6432 276
rect 6488 220 7492 276
rect 7548 220 7680 276
rect 7736 220 8740 276
rect 8796 220 8801 276
rect 6427 218 8801 220
rect 6427 215 6493 218
rect 7487 215 7553 218
rect 7675 215 7741 218
rect 8735 215 8801 218
rect 8923 278 8989 281
rect 9983 278 10049 281
rect 10171 278 10237 281
rect 11231 278 11297 281
rect 8923 276 11297 278
rect 8923 220 8928 276
rect 8984 220 9988 276
rect 10044 220 10176 276
rect 10232 220 11236 276
rect 11292 220 11297 276
rect 8923 218 11297 220
rect 8923 215 8989 218
rect 9983 215 10049 218
rect 10171 215 10237 218
rect 11231 215 11297 218
rect 11419 278 11485 281
rect 12479 278 12545 281
rect 12667 278 12733 281
rect 13727 278 13793 281
rect 11419 276 13793 278
rect 11419 220 11424 276
rect 11480 220 12484 276
rect 12540 220 12672 276
rect 12728 220 13732 276
rect 13788 220 13793 276
rect 11419 218 13793 220
rect 11419 215 11485 218
rect 12479 215 12545 218
rect 12667 215 12733 218
rect 13727 215 13793 218
rect 13915 278 13981 281
rect 14975 278 15041 281
rect 15163 278 15229 281
rect 16223 278 16289 281
rect 13915 276 16289 278
rect 13915 220 13920 276
rect 13976 220 14980 276
rect 15036 220 15168 276
rect 15224 220 16228 276
rect 16284 220 16289 276
rect 13915 218 16289 220
rect 13915 215 13981 218
rect 14975 215 15041 218
rect 15163 215 15229 218
rect 16223 215 16289 218
rect 16411 278 16477 281
rect 17471 278 17537 281
rect 17659 278 17725 281
rect 18719 278 18785 281
rect 16411 276 18785 278
rect 16411 220 16416 276
rect 16472 220 17476 276
rect 17532 220 17664 276
rect 17720 220 18724 276
rect 18780 220 18785 276
rect 16411 218 18785 220
rect 16411 215 16477 218
rect 17471 215 17537 218
rect 17659 215 17725 218
rect 18719 215 18785 218
rect 18907 278 18973 281
rect 19967 278 20033 281
rect 20155 278 20221 281
rect 21215 278 21281 281
rect 18907 276 21281 278
rect 18907 220 18912 276
rect 18968 220 19972 276
rect 20028 220 20160 276
rect 20216 220 21220 276
rect 21276 220 21281 276
rect 18907 218 21281 220
rect 18907 215 18973 218
rect 19967 215 20033 218
rect 20155 215 20221 218
rect 21215 215 21281 218
rect 21403 278 21469 281
rect 22463 278 22529 281
rect 22651 278 22717 281
rect 23711 278 23777 281
rect 21403 276 23777 278
rect 21403 220 21408 276
rect 21464 220 22468 276
rect 22524 220 22656 276
rect 22712 220 23716 276
rect 23772 220 23777 276
rect 21403 218 23777 220
rect 21403 215 21469 218
rect 22463 215 22529 218
rect 22651 215 22717 218
rect 23711 215 23777 218
rect 23899 278 23965 281
rect 24959 278 25025 281
rect 25147 278 25213 281
rect 26207 278 26273 281
rect 23899 276 26273 278
rect 23899 220 23904 276
rect 23960 220 24964 276
rect 25020 220 25152 276
rect 25208 220 26212 276
rect 26268 220 26273 276
rect 23899 218 26273 220
rect 23899 215 23965 218
rect 24959 215 25025 218
rect 25147 215 25213 218
rect 26207 215 26273 218
rect 26395 278 26461 281
rect 27455 278 27521 281
rect 27643 278 27709 281
rect 28703 278 28769 281
rect 26395 276 28769 278
rect 26395 220 26400 276
rect 26456 220 27460 276
rect 27516 220 27648 276
rect 27704 220 28708 276
rect 28764 220 28769 276
rect 26395 218 28769 220
rect 26395 215 26461 218
rect 27455 215 27521 218
rect 27643 215 27709 218
rect 28703 215 28769 218
rect 28891 278 28957 281
rect 29951 278 30017 281
rect 30139 278 30205 281
rect 31199 278 31265 281
rect 28891 276 31265 278
rect 28891 220 28896 276
rect 28952 220 29956 276
rect 30012 220 30144 276
rect 30200 220 31204 276
rect 31260 220 31265 276
rect 28891 218 31265 220
rect 28891 215 28957 218
rect 29951 215 30017 218
rect 30139 215 30205 218
rect 31199 215 31265 218
rect 31387 278 31453 281
rect 32447 278 32513 281
rect 32635 278 32701 281
rect 33695 278 33761 281
rect 31387 276 33761 278
rect 31387 220 31392 276
rect 31448 220 32452 276
rect 32508 220 32640 276
rect 32696 220 33700 276
rect 33756 220 33761 276
rect 31387 218 33761 220
rect 31387 215 31453 218
rect 32447 215 32513 218
rect 32635 215 32701 218
rect 33695 215 33761 218
rect 33883 278 33949 281
rect 34943 278 35009 281
rect 35131 278 35197 281
rect 36191 278 36257 281
rect 33883 276 36257 278
rect 33883 220 33888 276
rect 33944 220 34948 276
rect 35004 220 35136 276
rect 35192 220 36196 276
rect 36252 220 36257 276
rect 33883 218 36257 220
rect 33883 215 33949 218
rect 34943 215 35009 218
rect 35131 215 35197 218
rect 36191 215 36257 218
rect 36379 278 36445 281
rect 37439 278 37505 281
rect 37627 278 37693 281
rect 38687 278 38753 281
rect 36379 276 38753 278
rect 36379 220 36384 276
rect 36440 220 37444 276
rect 37500 220 37632 276
rect 37688 220 38692 276
rect 38748 220 38753 276
rect 36379 218 38753 220
rect 36379 215 36445 218
rect 37439 215 37505 218
rect 37627 215 37693 218
rect 38687 215 38753 218
rect 38875 278 38941 281
rect 39935 278 40001 281
rect 40123 278 40189 281
rect 41183 278 41249 281
rect 38875 276 41249 278
rect 38875 220 38880 276
rect 38936 220 39940 276
rect 39996 220 40128 276
rect 40184 220 41188 276
rect 41244 220 41249 276
rect 38875 218 41249 220
rect 38875 215 38941 218
rect 39935 215 40001 218
rect 40123 215 40189 218
rect 41183 215 41249 218
rect 41371 278 41437 281
rect 42431 278 42497 281
rect 42619 278 42685 281
rect 43679 278 43745 281
rect 41371 276 43745 278
rect 41371 220 41376 276
rect 41432 220 42436 276
rect 42492 220 42624 276
rect 42680 220 43684 276
rect 43740 220 43745 276
rect 41371 218 43745 220
rect 41371 215 41437 218
rect 42431 215 42497 218
rect 42619 215 42685 218
rect 43679 215 43745 218
rect 43867 278 43933 281
rect 44927 278 44993 281
rect 45115 278 45181 281
rect 46175 278 46241 281
rect 43867 276 46241 278
rect 43867 220 43872 276
rect 43928 220 44932 276
rect 44988 220 45120 276
rect 45176 220 46180 276
rect 46236 220 46241 276
rect 43867 218 46241 220
rect 43867 215 43933 218
rect 44927 215 44993 218
rect 45115 215 45181 218
rect 46175 215 46241 218
rect 46363 278 46429 281
rect 47423 278 47489 281
rect 47611 278 47677 281
rect 48671 278 48737 281
rect 46363 276 48737 278
rect 46363 220 46368 276
rect 46424 220 47428 276
rect 47484 220 47616 276
rect 47672 220 48676 276
rect 48732 220 48737 276
rect 46363 218 48737 220
rect 46363 215 46429 218
rect 47423 215 47489 218
rect 47611 215 47677 218
rect 48671 215 48737 218
rect 48859 278 48925 281
rect 49919 278 49985 281
rect 50107 278 50173 281
rect 51167 278 51233 281
rect 48859 276 51233 278
rect 48859 220 48864 276
rect 48920 220 49924 276
rect 49980 220 50112 276
rect 50168 220 51172 276
rect 51228 220 51233 276
rect 48859 218 51233 220
rect 48859 215 48925 218
rect 49919 215 49985 218
rect 50107 215 50173 218
rect 51167 215 51233 218
rect 51355 278 51421 281
rect 52415 278 52481 281
rect 52603 278 52669 281
rect 53663 278 53729 281
rect 51355 276 53729 278
rect 51355 220 51360 276
rect 51416 220 52420 276
rect 52476 220 52608 276
rect 52664 220 53668 276
rect 53724 220 53729 276
rect 51355 218 53729 220
rect 51355 215 51421 218
rect 52415 215 52481 218
rect 52603 215 52669 218
rect 53663 215 53729 218
rect 53851 278 53917 281
rect 54911 278 54977 281
rect 55099 278 55165 281
rect 56159 278 56225 281
rect 53851 276 56225 278
rect 53851 220 53856 276
rect 53912 220 54916 276
rect 54972 220 55104 276
rect 55160 220 56164 276
rect 56220 220 56225 276
rect 53851 218 56225 220
rect 53851 215 53917 218
rect 54911 215 54977 218
rect 55099 215 55165 218
rect 56159 215 56225 218
rect 56347 278 56413 281
rect 57407 278 57473 281
rect 57595 278 57661 281
rect 58655 278 58721 281
rect 56347 276 58721 278
rect 56347 220 56352 276
rect 56408 220 57412 276
rect 57468 220 57600 276
rect 57656 220 58660 276
rect 58716 220 58721 276
rect 56347 218 58721 220
rect 56347 215 56413 218
rect 57407 215 57473 218
rect 57595 215 57661 218
rect 58655 215 58721 218
rect 58843 278 58909 281
rect 59903 278 59969 281
rect 60091 278 60157 281
rect 61151 278 61217 281
rect 58843 276 61217 278
rect 58843 220 58848 276
rect 58904 220 59908 276
rect 59964 220 60096 276
rect 60152 220 61156 276
rect 61212 220 61217 276
rect 58843 218 61217 220
rect 58843 215 58909 218
rect 59903 215 59969 218
rect 60091 215 60157 218
rect 61151 215 61217 218
rect 61339 278 61405 281
rect 62399 278 62465 281
rect 62587 278 62653 281
rect 63647 278 63713 281
rect 61339 276 63713 278
rect 61339 220 61344 276
rect 61400 220 62404 276
rect 62460 220 62592 276
rect 62648 220 63652 276
rect 63708 220 63713 276
rect 61339 218 63713 220
rect 61339 215 61405 218
rect 62399 215 62465 218
rect 62587 215 62653 218
rect 63647 215 63713 218
rect 63835 278 63901 281
rect 64895 278 64961 281
rect 65083 278 65149 281
rect 66143 278 66209 281
rect 63835 276 66209 278
rect 63835 220 63840 276
rect 63896 220 64900 276
rect 64956 220 65088 276
rect 65144 220 66148 276
rect 66204 220 66209 276
rect 63835 218 66209 220
rect 63835 215 63901 218
rect 64895 215 64961 218
rect 65083 215 65149 218
rect 66143 215 66209 218
rect 66331 278 66397 281
rect 67391 278 67457 281
rect 67579 278 67645 281
rect 68639 278 68705 281
rect 66331 276 68705 278
rect 66331 220 66336 276
rect 66392 220 67396 276
rect 67452 220 67584 276
rect 67640 220 68644 276
rect 68700 220 68705 276
rect 66331 218 68705 220
rect 66331 215 66397 218
rect 67391 215 67457 218
rect 67579 215 67645 218
rect 68639 215 68705 218
rect 68827 278 68893 281
rect 69887 278 69953 281
rect 70075 278 70141 281
rect 71135 278 71201 281
rect 68827 276 71201 278
rect 68827 220 68832 276
rect 68888 220 69892 276
rect 69948 220 70080 276
rect 70136 220 71140 276
rect 71196 220 71201 276
rect 68827 218 71201 220
rect 68827 215 68893 218
rect 69887 215 69953 218
rect 70075 215 70141 218
rect 71135 215 71201 218
rect 71323 278 71389 281
rect 72383 278 72449 281
rect 72571 278 72637 281
rect 73631 278 73697 281
rect 71323 276 73697 278
rect 71323 220 71328 276
rect 71384 220 72388 276
rect 72444 220 72576 276
rect 72632 220 73636 276
rect 73692 220 73697 276
rect 71323 218 73697 220
rect 71323 215 71389 218
rect 72383 215 72449 218
rect 72571 215 72637 218
rect 73631 215 73697 218
rect 73819 278 73885 281
rect 74879 278 74945 281
rect 75067 278 75133 281
rect 76127 278 76193 281
rect 73819 276 76193 278
rect 73819 220 73824 276
rect 73880 220 74884 276
rect 74940 220 75072 276
rect 75128 220 76132 276
rect 76188 220 76193 276
rect 73819 218 76193 220
rect 73819 215 73885 218
rect 74879 215 74945 218
rect 75067 215 75133 218
rect 76127 215 76193 218
rect 76315 278 76381 281
rect 77375 278 77441 281
rect 77563 278 77629 281
rect 78623 278 78689 281
rect 76315 276 78689 278
rect 76315 220 76320 276
rect 76376 220 77380 276
rect 77436 220 77568 276
rect 77624 220 78628 276
rect 78684 220 78689 276
rect 76315 218 78689 220
rect 76315 215 76381 218
rect 77375 215 77441 218
rect 77563 215 77629 218
rect 78623 215 78689 218
rect 78811 278 78877 281
rect 79871 278 79937 281
rect 80059 278 80125 281
rect 81119 278 81185 281
rect 78811 276 81185 278
rect 78811 220 78816 276
rect 78872 220 79876 276
rect 79932 220 80064 276
rect 80120 220 81124 276
rect 81180 220 81185 276
rect 78811 218 81185 220
rect 78811 215 78877 218
rect 79871 215 79937 218
rect 80059 215 80125 218
rect 81119 215 81185 218
rect 1899 154 1965 157
rect 2031 154 2097 157
rect 3147 154 3213 157
rect 3279 154 3345 157
rect 1899 152 3345 154
rect 1899 96 1904 152
rect 1960 96 2036 152
rect 2092 96 3152 152
rect 3208 96 3284 152
rect 3340 96 3345 152
rect 1899 94 3345 96
rect 1899 91 1965 94
rect 2031 91 2097 94
rect 3147 91 3213 94
rect 3279 91 3345 94
rect 4395 154 4461 157
rect 4527 154 4593 157
rect 5643 154 5709 157
rect 5775 154 5841 157
rect 4395 152 5841 154
rect 4395 96 4400 152
rect 4456 96 4532 152
rect 4588 96 5648 152
rect 5704 96 5780 152
rect 5836 96 5841 152
rect 4395 94 5841 96
rect 4395 91 4461 94
rect 4527 91 4593 94
rect 5643 91 5709 94
rect 5775 91 5841 94
rect 6891 154 6957 157
rect 7023 154 7089 157
rect 8139 154 8205 157
rect 8271 154 8337 157
rect 6891 152 8337 154
rect 6891 96 6896 152
rect 6952 96 7028 152
rect 7084 96 8144 152
rect 8200 96 8276 152
rect 8332 96 8337 152
rect 6891 94 8337 96
rect 6891 91 6957 94
rect 7023 91 7089 94
rect 8139 91 8205 94
rect 8271 91 8337 94
rect 9387 154 9453 157
rect 9519 154 9585 157
rect 10635 154 10701 157
rect 10767 154 10833 157
rect 9387 152 10833 154
rect 9387 96 9392 152
rect 9448 96 9524 152
rect 9580 96 10640 152
rect 10696 96 10772 152
rect 10828 96 10833 152
rect 9387 94 10833 96
rect 9387 91 9453 94
rect 9519 91 9585 94
rect 10635 91 10701 94
rect 10767 91 10833 94
rect 11883 154 11949 157
rect 12015 154 12081 157
rect 13131 154 13197 157
rect 13263 154 13329 157
rect 11883 152 13329 154
rect 11883 96 11888 152
rect 11944 96 12020 152
rect 12076 96 13136 152
rect 13192 96 13268 152
rect 13324 96 13329 152
rect 11883 94 13329 96
rect 11883 91 11949 94
rect 12015 91 12081 94
rect 13131 91 13197 94
rect 13263 91 13329 94
rect 14379 154 14445 157
rect 14511 154 14577 157
rect 15627 154 15693 157
rect 15759 154 15825 157
rect 14379 152 15825 154
rect 14379 96 14384 152
rect 14440 96 14516 152
rect 14572 96 15632 152
rect 15688 96 15764 152
rect 15820 96 15825 152
rect 14379 94 15825 96
rect 14379 91 14445 94
rect 14511 91 14577 94
rect 15627 91 15693 94
rect 15759 91 15825 94
rect 16875 154 16941 157
rect 17007 154 17073 157
rect 18123 154 18189 157
rect 18255 154 18321 157
rect 16875 152 18321 154
rect 16875 96 16880 152
rect 16936 96 17012 152
rect 17068 96 18128 152
rect 18184 96 18260 152
rect 18316 96 18321 152
rect 16875 94 18321 96
rect 16875 91 16941 94
rect 17007 91 17073 94
rect 18123 91 18189 94
rect 18255 91 18321 94
rect 19371 154 19437 157
rect 19503 154 19569 157
rect 20619 154 20685 157
rect 20751 154 20817 157
rect 19371 152 20817 154
rect 19371 96 19376 152
rect 19432 96 19508 152
rect 19564 96 20624 152
rect 20680 96 20756 152
rect 20812 96 20817 152
rect 19371 94 20817 96
rect 19371 91 19437 94
rect 19503 91 19569 94
rect 20619 91 20685 94
rect 20751 91 20817 94
rect 21867 154 21933 157
rect 21999 154 22065 157
rect 23115 154 23181 157
rect 23247 154 23313 157
rect 21867 152 23313 154
rect 21867 96 21872 152
rect 21928 96 22004 152
rect 22060 96 23120 152
rect 23176 96 23252 152
rect 23308 96 23313 152
rect 21867 94 23313 96
rect 21867 91 21933 94
rect 21999 91 22065 94
rect 23115 91 23181 94
rect 23247 91 23313 94
rect 24363 154 24429 157
rect 24495 154 24561 157
rect 25611 154 25677 157
rect 25743 154 25809 157
rect 24363 152 25809 154
rect 24363 96 24368 152
rect 24424 96 24500 152
rect 24556 96 25616 152
rect 25672 96 25748 152
rect 25804 96 25809 152
rect 24363 94 25809 96
rect 24363 91 24429 94
rect 24495 91 24561 94
rect 25611 91 25677 94
rect 25743 91 25809 94
rect 26859 154 26925 157
rect 26991 154 27057 157
rect 28107 154 28173 157
rect 28239 154 28305 157
rect 26859 152 28305 154
rect 26859 96 26864 152
rect 26920 96 26996 152
rect 27052 96 28112 152
rect 28168 96 28244 152
rect 28300 96 28305 152
rect 26859 94 28305 96
rect 26859 91 26925 94
rect 26991 91 27057 94
rect 28107 91 28173 94
rect 28239 91 28305 94
rect 29355 154 29421 157
rect 29487 154 29553 157
rect 30603 154 30669 157
rect 30735 154 30801 157
rect 29355 152 30801 154
rect 29355 96 29360 152
rect 29416 96 29492 152
rect 29548 96 30608 152
rect 30664 96 30740 152
rect 30796 96 30801 152
rect 29355 94 30801 96
rect 29355 91 29421 94
rect 29487 91 29553 94
rect 30603 91 30669 94
rect 30735 91 30801 94
rect 31851 154 31917 157
rect 31983 154 32049 157
rect 33099 154 33165 157
rect 33231 154 33297 157
rect 31851 152 33297 154
rect 31851 96 31856 152
rect 31912 96 31988 152
rect 32044 96 33104 152
rect 33160 96 33236 152
rect 33292 96 33297 152
rect 31851 94 33297 96
rect 31851 91 31917 94
rect 31983 91 32049 94
rect 33099 91 33165 94
rect 33231 91 33297 94
rect 34347 154 34413 157
rect 34479 154 34545 157
rect 35595 154 35661 157
rect 35727 154 35793 157
rect 34347 152 35793 154
rect 34347 96 34352 152
rect 34408 96 34484 152
rect 34540 96 35600 152
rect 35656 96 35732 152
rect 35788 96 35793 152
rect 34347 94 35793 96
rect 34347 91 34413 94
rect 34479 91 34545 94
rect 35595 91 35661 94
rect 35727 91 35793 94
rect 36843 154 36909 157
rect 36975 154 37041 157
rect 38091 154 38157 157
rect 38223 154 38289 157
rect 36843 152 38289 154
rect 36843 96 36848 152
rect 36904 96 36980 152
rect 37036 96 38096 152
rect 38152 96 38228 152
rect 38284 96 38289 152
rect 36843 94 38289 96
rect 36843 91 36909 94
rect 36975 91 37041 94
rect 38091 91 38157 94
rect 38223 91 38289 94
rect 39339 154 39405 157
rect 39471 154 39537 157
rect 40587 154 40653 157
rect 40719 154 40785 157
rect 39339 152 40785 154
rect 39339 96 39344 152
rect 39400 96 39476 152
rect 39532 96 40592 152
rect 40648 96 40724 152
rect 40780 96 40785 152
rect 39339 94 40785 96
rect 39339 91 39405 94
rect 39471 91 39537 94
rect 40587 91 40653 94
rect 40719 91 40785 94
rect 41835 154 41901 157
rect 41967 154 42033 157
rect 43083 154 43149 157
rect 43215 154 43281 157
rect 41835 152 43281 154
rect 41835 96 41840 152
rect 41896 96 41972 152
rect 42028 96 43088 152
rect 43144 96 43220 152
rect 43276 96 43281 152
rect 41835 94 43281 96
rect 41835 91 41901 94
rect 41967 91 42033 94
rect 43083 91 43149 94
rect 43215 91 43281 94
rect 44331 154 44397 157
rect 44463 154 44529 157
rect 45579 154 45645 157
rect 45711 154 45777 157
rect 44331 152 45777 154
rect 44331 96 44336 152
rect 44392 96 44468 152
rect 44524 96 45584 152
rect 45640 96 45716 152
rect 45772 96 45777 152
rect 44331 94 45777 96
rect 44331 91 44397 94
rect 44463 91 44529 94
rect 45579 91 45645 94
rect 45711 91 45777 94
rect 46827 154 46893 157
rect 46959 154 47025 157
rect 48075 154 48141 157
rect 48207 154 48273 157
rect 46827 152 48273 154
rect 46827 96 46832 152
rect 46888 96 46964 152
rect 47020 96 48080 152
rect 48136 96 48212 152
rect 48268 96 48273 152
rect 46827 94 48273 96
rect 46827 91 46893 94
rect 46959 91 47025 94
rect 48075 91 48141 94
rect 48207 91 48273 94
rect 49323 154 49389 157
rect 49455 154 49521 157
rect 50571 154 50637 157
rect 50703 154 50769 157
rect 49323 152 50769 154
rect 49323 96 49328 152
rect 49384 96 49460 152
rect 49516 96 50576 152
rect 50632 96 50708 152
rect 50764 96 50769 152
rect 49323 94 50769 96
rect 49323 91 49389 94
rect 49455 91 49521 94
rect 50571 91 50637 94
rect 50703 91 50769 94
rect 51819 154 51885 157
rect 51951 154 52017 157
rect 53067 154 53133 157
rect 53199 154 53265 157
rect 51819 152 53265 154
rect 51819 96 51824 152
rect 51880 96 51956 152
rect 52012 96 53072 152
rect 53128 96 53204 152
rect 53260 96 53265 152
rect 51819 94 53265 96
rect 51819 91 51885 94
rect 51951 91 52017 94
rect 53067 91 53133 94
rect 53199 91 53265 94
rect 54315 154 54381 157
rect 54447 154 54513 157
rect 55563 154 55629 157
rect 55695 154 55761 157
rect 54315 152 55761 154
rect 54315 96 54320 152
rect 54376 96 54452 152
rect 54508 96 55568 152
rect 55624 96 55700 152
rect 55756 96 55761 152
rect 54315 94 55761 96
rect 54315 91 54381 94
rect 54447 91 54513 94
rect 55563 91 55629 94
rect 55695 91 55761 94
rect 56811 154 56877 157
rect 56943 154 57009 157
rect 58059 154 58125 157
rect 58191 154 58257 157
rect 56811 152 58257 154
rect 56811 96 56816 152
rect 56872 96 56948 152
rect 57004 96 58064 152
rect 58120 96 58196 152
rect 58252 96 58257 152
rect 56811 94 58257 96
rect 56811 91 56877 94
rect 56943 91 57009 94
rect 58059 91 58125 94
rect 58191 91 58257 94
rect 59307 154 59373 157
rect 59439 154 59505 157
rect 60555 154 60621 157
rect 60687 154 60753 157
rect 59307 152 60753 154
rect 59307 96 59312 152
rect 59368 96 59444 152
rect 59500 96 60560 152
rect 60616 96 60692 152
rect 60748 96 60753 152
rect 59307 94 60753 96
rect 59307 91 59373 94
rect 59439 91 59505 94
rect 60555 91 60621 94
rect 60687 91 60753 94
rect 61803 154 61869 157
rect 61935 154 62001 157
rect 63051 154 63117 157
rect 63183 154 63249 157
rect 61803 152 63249 154
rect 61803 96 61808 152
rect 61864 96 61940 152
rect 61996 96 63056 152
rect 63112 96 63188 152
rect 63244 96 63249 152
rect 61803 94 63249 96
rect 61803 91 61869 94
rect 61935 91 62001 94
rect 63051 91 63117 94
rect 63183 91 63249 94
rect 64299 154 64365 157
rect 64431 154 64497 157
rect 65547 154 65613 157
rect 65679 154 65745 157
rect 64299 152 65745 154
rect 64299 96 64304 152
rect 64360 96 64436 152
rect 64492 96 65552 152
rect 65608 96 65684 152
rect 65740 96 65745 152
rect 64299 94 65745 96
rect 64299 91 64365 94
rect 64431 91 64497 94
rect 65547 91 65613 94
rect 65679 91 65745 94
rect 66795 154 66861 157
rect 66927 154 66993 157
rect 68043 154 68109 157
rect 68175 154 68241 157
rect 66795 152 68241 154
rect 66795 96 66800 152
rect 66856 96 66932 152
rect 66988 96 68048 152
rect 68104 96 68180 152
rect 68236 96 68241 152
rect 66795 94 68241 96
rect 66795 91 66861 94
rect 66927 91 66993 94
rect 68043 91 68109 94
rect 68175 91 68241 94
rect 69291 154 69357 157
rect 69423 154 69489 157
rect 70539 154 70605 157
rect 70671 154 70737 157
rect 69291 152 70737 154
rect 69291 96 69296 152
rect 69352 96 69428 152
rect 69484 96 70544 152
rect 70600 96 70676 152
rect 70732 96 70737 152
rect 69291 94 70737 96
rect 69291 91 69357 94
rect 69423 91 69489 94
rect 70539 91 70605 94
rect 70671 91 70737 94
rect 71787 154 71853 157
rect 71919 154 71985 157
rect 73035 154 73101 157
rect 73167 154 73233 157
rect 71787 152 73233 154
rect 71787 96 71792 152
rect 71848 96 71924 152
rect 71980 96 73040 152
rect 73096 96 73172 152
rect 73228 96 73233 152
rect 71787 94 73233 96
rect 71787 91 71853 94
rect 71919 91 71985 94
rect 73035 91 73101 94
rect 73167 91 73233 94
rect 74283 154 74349 157
rect 74415 154 74481 157
rect 75531 154 75597 157
rect 75663 154 75729 157
rect 74283 152 75729 154
rect 74283 96 74288 152
rect 74344 96 74420 152
rect 74476 96 75536 152
rect 75592 96 75668 152
rect 75724 96 75729 152
rect 74283 94 75729 96
rect 74283 91 74349 94
rect 74415 91 74481 94
rect 75531 91 75597 94
rect 75663 91 75729 94
rect 76779 154 76845 157
rect 76911 154 76977 157
rect 78027 154 78093 157
rect 78159 154 78225 157
rect 76779 152 78225 154
rect 76779 96 76784 152
rect 76840 96 76916 152
rect 76972 96 78032 152
rect 78088 96 78164 152
rect 78220 96 78225 152
rect 76779 94 78225 96
rect 76779 91 76845 94
rect 76911 91 76977 94
rect 78027 91 78093 94
rect 78159 91 78225 94
rect 79275 154 79341 157
rect 79407 154 79473 157
rect 80523 154 80589 157
rect 80655 154 80721 157
rect 79275 152 80721 154
rect 79275 96 79280 152
rect 79336 96 79412 152
rect 79468 96 80528 152
rect 80584 96 80660 152
rect 80716 96 80721 152
rect 79275 94 80721 96
rect 79275 91 79341 94
rect 79407 91 79473 94
rect 80523 91 80589 94
rect 80655 91 80721 94
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_0
timestamp 1676037725
transform -1 0 6366 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_1
timestamp 1676037725
transform 1 0 5118 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_2
timestamp 1676037725
transform -1 0 5118 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_3
timestamp 1676037725
transform 1 0 3870 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_4
timestamp 1676037725
transform -1 0 3870 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_5
timestamp 1676037725
transform 1 0 2622 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_6
timestamp 1676037725
transform -1 0 2622 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_7
timestamp 1676037725
transform 1 0 1374 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_8
timestamp 1676037725
transform -1 0 11358 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_9
timestamp 1676037725
transform 1 0 10110 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_10
timestamp 1676037725
transform -1 0 10110 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_11
timestamp 1676037725
transform 1 0 8862 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_12
timestamp 1676037725
transform -1 0 8862 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_13
timestamp 1676037725
transform 1 0 7614 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_14
timestamp 1676037725
transform -1 0 7614 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_15
timestamp 1676037725
transform 1 0 6366 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_16
timestamp 1676037725
transform -1 0 16350 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_17
timestamp 1676037725
transform 1 0 15102 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_18
timestamp 1676037725
transform -1 0 15102 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_19
timestamp 1676037725
transform 1 0 13854 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_20
timestamp 1676037725
transform -1 0 13854 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_21
timestamp 1676037725
transform 1 0 12606 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_22
timestamp 1676037725
transform -1 0 12606 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_23
timestamp 1676037725
transform 1 0 11358 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_24
timestamp 1676037725
transform -1 0 21342 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_25
timestamp 1676037725
transform 1 0 20094 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_26
timestamp 1676037725
transform -1 0 20094 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_27
timestamp 1676037725
transform 1 0 18846 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_28
timestamp 1676037725
transform -1 0 18846 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_29
timestamp 1676037725
transform 1 0 17598 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_30
timestamp 1676037725
transform -1 0 17598 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_31
timestamp 1676037725
transform 1 0 16350 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_32
timestamp 1676037725
transform -1 0 26334 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_33
timestamp 1676037725
transform 1 0 25086 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_34
timestamp 1676037725
transform -1 0 25086 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_35
timestamp 1676037725
transform 1 0 23838 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_36
timestamp 1676037725
transform -1 0 23838 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_37
timestamp 1676037725
transform 1 0 22590 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_38
timestamp 1676037725
transform -1 0 22590 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_39
timestamp 1676037725
transform 1 0 21342 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_40
timestamp 1676037725
transform -1 0 31326 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_41
timestamp 1676037725
transform 1 0 30078 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_42
timestamp 1676037725
transform -1 0 30078 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_43
timestamp 1676037725
transform 1 0 28830 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_44
timestamp 1676037725
transform -1 0 28830 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_45
timestamp 1676037725
transform 1 0 27582 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_46
timestamp 1676037725
transform -1 0 27582 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_47
timestamp 1676037725
transform 1 0 26334 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_48
timestamp 1676037725
transform -1 0 36318 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_49
timestamp 1676037725
transform 1 0 35070 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_50
timestamp 1676037725
transform -1 0 35070 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_51
timestamp 1676037725
transform 1 0 33822 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_52
timestamp 1676037725
transform -1 0 33822 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_53
timestamp 1676037725
transform 1 0 32574 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_54
timestamp 1676037725
transform -1 0 32574 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_55
timestamp 1676037725
transform 1 0 31326 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_56
timestamp 1676037725
transform -1 0 41310 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_57
timestamp 1676037725
transform 1 0 40062 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_58
timestamp 1676037725
transform -1 0 40062 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_59
timestamp 1676037725
transform 1 0 38814 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_60
timestamp 1676037725
transform -1 0 38814 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_61
timestamp 1676037725
transform 1 0 37566 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_62
timestamp 1676037725
transform -1 0 37566 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_63
timestamp 1676037725
transform 1 0 36318 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_64
timestamp 1676037725
transform -1 0 46302 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_65
timestamp 1676037725
transform 1 0 45054 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_66
timestamp 1676037725
transform -1 0 45054 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_67
timestamp 1676037725
transform 1 0 43806 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_68
timestamp 1676037725
transform -1 0 43806 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_69
timestamp 1676037725
transform 1 0 42558 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_70
timestamp 1676037725
transform -1 0 42558 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_71
timestamp 1676037725
transform 1 0 41310 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_72
timestamp 1676037725
transform -1 0 51294 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_73
timestamp 1676037725
transform 1 0 50046 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_74
timestamp 1676037725
transform -1 0 50046 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_75
timestamp 1676037725
transform 1 0 48798 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_76
timestamp 1676037725
transform -1 0 48798 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_77
timestamp 1676037725
transform 1 0 47550 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_78
timestamp 1676037725
transform -1 0 47550 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_79
timestamp 1676037725
transform 1 0 46302 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_80
timestamp 1676037725
transform -1 0 56286 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_81
timestamp 1676037725
transform 1 0 55038 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_82
timestamp 1676037725
transform -1 0 55038 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_83
timestamp 1676037725
transform 1 0 53790 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_84
timestamp 1676037725
transform -1 0 53790 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_85
timestamp 1676037725
transform 1 0 52542 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_86
timestamp 1676037725
transform -1 0 52542 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_87
timestamp 1676037725
transform 1 0 51294 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_88
timestamp 1676037725
transform -1 0 61278 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_89
timestamp 1676037725
transform 1 0 60030 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_90
timestamp 1676037725
transform -1 0 60030 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_91
timestamp 1676037725
transform 1 0 58782 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_92
timestamp 1676037725
transform -1 0 58782 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_93
timestamp 1676037725
transform 1 0 57534 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_94
timestamp 1676037725
transform -1 0 57534 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_95
timestamp 1676037725
transform 1 0 56286 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_96
timestamp 1676037725
transform -1 0 66270 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_97
timestamp 1676037725
transform 1 0 65022 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_98
timestamp 1676037725
transform -1 0 65022 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_99
timestamp 1676037725
transform 1 0 63774 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_100
timestamp 1676037725
transform -1 0 63774 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_101
timestamp 1676037725
transform 1 0 62526 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_102
timestamp 1676037725
transform -1 0 62526 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_103
timestamp 1676037725
transform 1 0 61278 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_104
timestamp 1676037725
transform -1 0 71262 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_105
timestamp 1676037725
transform 1 0 70014 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_106
timestamp 1676037725
transform -1 0 70014 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_107
timestamp 1676037725
transform 1 0 68766 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_108
timestamp 1676037725
transform -1 0 68766 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_109
timestamp 1676037725
transform 1 0 67518 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_110
timestamp 1676037725
transform -1 0 67518 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_111
timestamp 1676037725
transform 1 0 66270 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_112
timestamp 1676037725
transform -1 0 76254 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_113
timestamp 1676037725
transform 1 0 75006 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_114
timestamp 1676037725
transform -1 0 75006 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_115
timestamp 1676037725
transform 1 0 73758 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_116
timestamp 1676037725
transform -1 0 73758 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_117
timestamp 1676037725
transform 1 0 72510 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_118
timestamp 1676037725
transform -1 0 72510 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_119
timestamp 1676037725
transform 1 0 71262 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_120
timestamp 1676037725
transform -1 0 81246 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_121
timestamp 1676037725
transform 1 0 79998 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_122
timestamp 1676037725
transform -1 0 79998 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_123
timestamp 1676037725
transform 1 0 78750 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_124
timestamp 1676037725
transform -1 0 78750 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_125
timestamp 1676037725
transform 1 0 77502 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_126
timestamp 1676037725
transform -1 0 77502 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_127
timestamp 1676037725
transform 1 0 76254 0 1 868
box 65 0 675 1316
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_0
timestamp 1676037725
transform 1 0 4773 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_1
timestamp 1676037725
transform 1 0 4149 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_2
timestamp 1676037725
transform 1 0 3525 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_3
timestamp 1676037725
transform 1 0 2901 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_4
timestamp 1676037725
transform 1 0 2277 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_5
timestamp 1676037725
transform 1 0 1653 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_6
timestamp 1676037725
transform 1 0 6021 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_7
timestamp 1676037725
transform 1 0 5397 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_8
timestamp 1676037725
transform 1 0 11013 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_9
timestamp 1676037725
transform 1 0 10389 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_10
timestamp 1676037725
transform 1 0 9765 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_11
timestamp 1676037725
transform 1 0 9141 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_12
timestamp 1676037725
transform 1 0 8517 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_13
timestamp 1676037725
transform 1 0 7893 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_14
timestamp 1676037725
transform 1 0 7269 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_15
timestamp 1676037725
transform 1 0 6645 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_16
timestamp 1676037725
transform 1 0 16005 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_17
timestamp 1676037725
transform 1 0 15381 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_18
timestamp 1676037725
transform 1 0 14757 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_19
timestamp 1676037725
transform 1 0 14133 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_20
timestamp 1676037725
transform 1 0 13509 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_21
timestamp 1676037725
transform 1 0 12885 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_22
timestamp 1676037725
transform 1 0 12261 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_23
timestamp 1676037725
transform 1 0 11637 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_24
timestamp 1676037725
transform 1 0 20997 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_25
timestamp 1676037725
transform 1 0 20373 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_26
timestamp 1676037725
transform 1 0 19749 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_27
timestamp 1676037725
transform 1 0 19125 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_28
timestamp 1676037725
transform 1 0 18501 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_29
timestamp 1676037725
transform 1 0 17877 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_30
timestamp 1676037725
transform 1 0 17253 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_31
timestamp 1676037725
transform 1 0 16629 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_32
timestamp 1676037725
transform 1 0 23493 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_33
timestamp 1676037725
transform 1 0 22869 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_34
timestamp 1676037725
transform 1 0 22245 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_35
timestamp 1676037725
transform 1 0 21621 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_36
timestamp 1676037725
transform 1 0 25989 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_37
timestamp 1676037725
transform 1 0 25365 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_38
timestamp 1676037725
transform 1 0 24741 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_39
timestamp 1676037725
transform 1 0 24117 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_40
timestamp 1676037725
transform 1 0 30981 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_41
timestamp 1676037725
transform 1 0 30357 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_42
timestamp 1676037725
transform 1 0 29733 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_43
timestamp 1676037725
transform 1 0 29109 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_44
timestamp 1676037725
transform 1 0 28485 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_45
timestamp 1676037725
transform 1 0 27861 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_46
timestamp 1676037725
transform 1 0 27237 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_47
timestamp 1676037725
transform 1 0 26613 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_48
timestamp 1676037725
transform 1 0 32229 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_49
timestamp 1676037725
transform 1 0 31605 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_50
timestamp 1676037725
transform 1 0 35973 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_51
timestamp 1676037725
transform 1 0 35349 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_52
timestamp 1676037725
transform 1 0 34725 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_53
timestamp 1676037725
transform 1 0 34101 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_54
timestamp 1676037725
transform 1 0 33477 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_55
timestamp 1676037725
transform 1 0 32853 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_56
timestamp 1676037725
transform 1 0 40965 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_57
timestamp 1676037725
transform 1 0 40341 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_58
timestamp 1676037725
transform 1 0 39717 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_59
timestamp 1676037725
transform 1 0 39093 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_60
timestamp 1676037725
transform 1 0 38469 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_61
timestamp 1676037725
transform 1 0 37845 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_62
timestamp 1676037725
transform 1 0 37221 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_63
timestamp 1676037725
transform 1 0 36597 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_64
timestamp 1676037725
transform 1 0 45957 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_65
timestamp 1676037725
transform 1 0 45333 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_66
timestamp 1676037725
transform 1 0 44709 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_67
timestamp 1676037725
transform 1 0 44085 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_68
timestamp 1676037725
transform 1 0 43461 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_69
timestamp 1676037725
transform 1 0 42837 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_70
timestamp 1676037725
transform 1 0 42213 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_71
timestamp 1676037725
transform 1 0 41589 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_72
timestamp 1676037725
transform 1 0 50949 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_73
timestamp 1676037725
transform 1 0 50325 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_74
timestamp 1676037725
transform 1 0 49701 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_75
timestamp 1676037725
transform 1 0 49077 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_76
timestamp 1676037725
transform 1 0 48453 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_77
timestamp 1676037725
transform 1 0 47829 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_78
timestamp 1676037725
transform 1 0 47205 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_79
timestamp 1676037725
transform 1 0 46581 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_80
timestamp 1676037725
transform 1 0 52197 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_81
timestamp 1676037725
transform 1 0 51573 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_82
timestamp 1676037725
transform 1 0 55941 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_83
timestamp 1676037725
transform 1 0 55317 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_84
timestamp 1676037725
transform 1 0 54693 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_85
timestamp 1676037725
transform 1 0 54069 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_86
timestamp 1676037725
transform 1 0 53445 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_87
timestamp 1676037725
transform 1 0 52821 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_88
timestamp 1676037725
transform 1 0 60933 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_89
timestamp 1676037725
transform 1 0 60309 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_90
timestamp 1676037725
transform 1 0 59685 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_91
timestamp 1676037725
transform 1 0 59061 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_92
timestamp 1676037725
transform 1 0 58437 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_93
timestamp 1676037725
transform 1 0 57813 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_94
timestamp 1676037725
transform 1 0 57189 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_95
timestamp 1676037725
transform 1 0 56565 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_96
timestamp 1676037725
transform 1 0 65925 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_97
timestamp 1676037725
transform 1 0 65301 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_98
timestamp 1676037725
transform 1 0 64677 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_99
timestamp 1676037725
transform 1 0 64053 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_100
timestamp 1676037725
transform 1 0 63429 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_101
timestamp 1676037725
transform 1 0 62805 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_102
timestamp 1676037725
transform 1 0 62181 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_103
timestamp 1676037725
transform 1 0 61557 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_104
timestamp 1676037725
transform 1 0 70917 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_105
timestamp 1676037725
transform 1 0 70293 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_106
timestamp 1676037725
transform 1 0 69669 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_107
timestamp 1676037725
transform 1 0 69045 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_108
timestamp 1676037725
transform 1 0 68421 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_109
timestamp 1676037725
transform 1 0 67797 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_110
timestamp 1676037725
transform 1 0 67173 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_111
timestamp 1676037725
transform 1 0 66549 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_112
timestamp 1676037725
transform 1 0 73413 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_113
timestamp 1676037725
transform 1 0 72789 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_114
timestamp 1676037725
transform 1 0 72165 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_115
timestamp 1676037725
transform 1 0 71541 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_116
timestamp 1676037725
transform 1 0 75909 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_117
timestamp 1676037725
transform 1 0 75285 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_118
timestamp 1676037725
transform 1 0 74661 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_119
timestamp 1676037725
transform 1 0 74037 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_120
timestamp 1676037725
transform 1 0 80901 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_121
timestamp 1676037725
transform 1 0 80277 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_122
timestamp 1676037725
transform 1 0 79653 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_123
timestamp 1676037725
transform 1 0 79029 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_124
timestamp 1676037725
transform 1 0 78405 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_125
timestamp 1676037725
transform 1 0 77781 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_126
timestamp 1676037725
transform 1 0 77157 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_24  sky130_sram_2kbyte_1rw1r_32x512_8_contact_24_127
timestamp 1676037725
transform 1 0 76533 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_0
timestamp 1676037725
transform 1 0 4777 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_1
timestamp 1676037725
transform 1 0 4153 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_2
timestamp 1676037725
transform 1 0 3529 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_3
timestamp 1676037725
transform 1 0 2905 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_4
timestamp 1676037725
transform 1 0 2281 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_5
timestamp 1676037725
transform 1 0 1657 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_6
timestamp 1676037725
transform 1 0 6025 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_7
timestamp 1676037725
transform 1 0 5401 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_8
timestamp 1676037725
transform 1 0 11017 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_9
timestamp 1676037725
transform 1 0 10393 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_10
timestamp 1676037725
transform 1 0 9769 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_11
timestamp 1676037725
transform 1 0 9145 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_12
timestamp 1676037725
transform 1 0 8521 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_13
timestamp 1676037725
transform 1 0 7897 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_14
timestamp 1676037725
transform 1 0 7273 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_15
timestamp 1676037725
transform 1 0 6649 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_16
timestamp 1676037725
transform 1 0 16009 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_17
timestamp 1676037725
transform 1 0 15385 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_18
timestamp 1676037725
transform 1 0 14761 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_19
timestamp 1676037725
transform 1 0 14137 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_20
timestamp 1676037725
transform 1 0 13513 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_21
timestamp 1676037725
transform 1 0 12889 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_22
timestamp 1676037725
transform 1 0 12265 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_23
timestamp 1676037725
transform 1 0 11641 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_24
timestamp 1676037725
transform 1 0 21001 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_25
timestamp 1676037725
transform 1 0 20377 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_26
timestamp 1676037725
transform 1 0 19753 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_27
timestamp 1676037725
transform 1 0 19129 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_28
timestamp 1676037725
transform 1 0 18505 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_29
timestamp 1676037725
transform 1 0 17881 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_30
timestamp 1676037725
transform 1 0 17257 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_31
timestamp 1676037725
transform 1 0 16633 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_32
timestamp 1676037725
transform 1 0 23497 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_33
timestamp 1676037725
transform 1 0 22873 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_34
timestamp 1676037725
transform 1 0 22249 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_35
timestamp 1676037725
transform 1 0 21625 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_36
timestamp 1676037725
transform 1 0 25993 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_37
timestamp 1676037725
transform 1 0 25369 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_38
timestamp 1676037725
transform 1 0 24745 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_39
timestamp 1676037725
transform 1 0 24121 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_40
timestamp 1676037725
transform 1 0 30985 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_41
timestamp 1676037725
transform 1 0 30361 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_42
timestamp 1676037725
transform 1 0 29737 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_43
timestamp 1676037725
transform 1 0 29113 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_44
timestamp 1676037725
transform 1 0 28489 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_45
timestamp 1676037725
transform 1 0 27865 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_46
timestamp 1676037725
transform 1 0 27241 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_47
timestamp 1676037725
transform 1 0 26617 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_48
timestamp 1676037725
transform 1 0 32233 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_49
timestamp 1676037725
transform 1 0 31609 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_50
timestamp 1676037725
transform 1 0 35977 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_51
timestamp 1676037725
transform 1 0 35353 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_52
timestamp 1676037725
transform 1 0 34729 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_53
timestamp 1676037725
transform 1 0 34105 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_54
timestamp 1676037725
transform 1 0 33481 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_55
timestamp 1676037725
transform 1 0 32857 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_56
timestamp 1676037725
transform 1 0 40969 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_57
timestamp 1676037725
transform 1 0 40345 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_58
timestamp 1676037725
transform 1 0 39721 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_59
timestamp 1676037725
transform 1 0 39097 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_60
timestamp 1676037725
transform 1 0 38473 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_61
timestamp 1676037725
transform 1 0 37849 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_62
timestamp 1676037725
transform 1 0 37225 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_63
timestamp 1676037725
transform 1 0 36601 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_64
timestamp 1676037725
transform 1 0 45961 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_65
timestamp 1676037725
transform 1 0 45337 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_66
timestamp 1676037725
transform 1 0 44713 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_67
timestamp 1676037725
transform 1 0 44089 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_68
timestamp 1676037725
transform 1 0 43465 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_69
timestamp 1676037725
transform 1 0 42841 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_70
timestamp 1676037725
transform 1 0 42217 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_71
timestamp 1676037725
transform 1 0 41593 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_72
timestamp 1676037725
transform 1 0 50953 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_73
timestamp 1676037725
transform 1 0 50329 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_74
timestamp 1676037725
transform 1 0 49705 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_75
timestamp 1676037725
transform 1 0 49081 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_76
timestamp 1676037725
transform 1 0 48457 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_77
timestamp 1676037725
transform 1 0 47833 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_78
timestamp 1676037725
transform 1 0 47209 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_79
timestamp 1676037725
transform 1 0 46585 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_80
timestamp 1676037725
transform 1 0 52201 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_81
timestamp 1676037725
transform 1 0 51577 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_82
timestamp 1676037725
transform 1 0 55945 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_83
timestamp 1676037725
transform 1 0 55321 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_84
timestamp 1676037725
transform 1 0 54697 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_85
timestamp 1676037725
transform 1 0 54073 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_86
timestamp 1676037725
transform 1 0 53449 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_87
timestamp 1676037725
transform 1 0 52825 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_88
timestamp 1676037725
transform 1 0 60937 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_89
timestamp 1676037725
transform 1 0 60313 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_90
timestamp 1676037725
transform 1 0 59689 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_91
timestamp 1676037725
transform 1 0 59065 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_92
timestamp 1676037725
transform 1 0 58441 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_93
timestamp 1676037725
transform 1 0 57817 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_94
timestamp 1676037725
transform 1 0 57193 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_95
timestamp 1676037725
transform 1 0 56569 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_96
timestamp 1676037725
transform 1 0 65929 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_97
timestamp 1676037725
transform 1 0 65305 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_98
timestamp 1676037725
transform 1 0 64681 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_99
timestamp 1676037725
transform 1 0 64057 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_100
timestamp 1676037725
transform 1 0 63433 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_101
timestamp 1676037725
transform 1 0 62809 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_102
timestamp 1676037725
transform 1 0 62185 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_103
timestamp 1676037725
transform 1 0 61561 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_104
timestamp 1676037725
transform 1 0 70921 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_105
timestamp 1676037725
transform 1 0 70297 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_106
timestamp 1676037725
transform 1 0 69673 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_107
timestamp 1676037725
transform 1 0 69049 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_108
timestamp 1676037725
transform 1 0 68425 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_109
timestamp 1676037725
transform 1 0 67801 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_110
timestamp 1676037725
transform 1 0 67177 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_111
timestamp 1676037725
transform 1 0 66553 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_112
timestamp 1676037725
transform 1 0 73417 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_113
timestamp 1676037725
transform 1 0 72793 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_114
timestamp 1676037725
transform 1 0 72169 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_115
timestamp 1676037725
transform 1 0 71545 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_116
timestamp 1676037725
transform 1 0 75913 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_117
timestamp 1676037725
transform 1 0 75289 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_118
timestamp 1676037725
transform 1 0 74665 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_119
timestamp 1676037725
transform 1 0 74041 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_120
timestamp 1676037725
transform 1 0 80905 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_121
timestamp 1676037725
transform 1 0 80281 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_122
timestamp 1676037725
transform 1 0 79657 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_123
timestamp 1676037725
transform 1 0 79033 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_124
timestamp 1676037725
transform 1 0 78409 0 1 741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_125
timestamp 1676037725
transform 1 0 77785 0 1 617
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_126
timestamp 1676037725
transform 1 0 77161 0 1 493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_25  sky130_sram_2kbyte_1rw1r_32x512_8_contact_25_127
timestamp 1676037725
transform 1 0 76537 0 1 369
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_0
timestamp 1676037725
transform 1 0 5776 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_1
timestamp 1676037725
transform 1 0 6240 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_2
timestamp 1676037725
transform 1 0 5644 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_3
timestamp 1676037725
transform 1 0 5180 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_4
timestamp 1676037725
transform 1 0 4528 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_5
timestamp 1676037725
transform 1 0 4992 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_6
timestamp 1676037725
transform 1 0 4396 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_7
timestamp 1676037725
transform 1 0 3932 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_8
timestamp 1676037725
transform 1 0 3280 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_9
timestamp 1676037725
transform 1 0 3744 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_10
timestamp 1676037725
transform 1 0 3148 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_11
timestamp 1676037725
transform 1 0 2684 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_12
timestamp 1676037725
transform 1 0 2032 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_13
timestamp 1676037725
transform 1 0 2496 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_14
timestamp 1676037725
transform 1 0 1900 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_15
timestamp 1676037725
transform 1 0 1436 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_16
timestamp 1676037725
transform 1 0 4774 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_17
timestamp 1676037725
transform 1 0 4150 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_18
timestamp 1676037725
transform 1 0 3526 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_19
timestamp 1676037725
transform 1 0 2902 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_20
timestamp 1676037725
transform 1 0 2278 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_21
timestamp 1676037725
transform 1 0 1654 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_22
timestamp 1676037725
transform 1 0 6022 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_23
timestamp 1676037725
transform 1 0 5398 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_24
timestamp 1676037725
transform 1 0 10768 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_25
timestamp 1676037725
transform 1 0 11232 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_26
timestamp 1676037725
transform 1 0 10636 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_27
timestamp 1676037725
transform 1 0 10172 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_28
timestamp 1676037725
transform 1 0 9520 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_29
timestamp 1676037725
transform 1 0 9984 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_30
timestamp 1676037725
transform 1 0 9388 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_31
timestamp 1676037725
transform 1 0 8924 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_32
timestamp 1676037725
transform 1 0 11014 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_33
timestamp 1676037725
transform 1 0 10390 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_34
timestamp 1676037725
transform 1 0 9766 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_35
timestamp 1676037725
transform 1 0 9142 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_36
timestamp 1676037725
transform 1 0 8518 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_37
timestamp 1676037725
transform 1 0 7894 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_38
timestamp 1676037725
transform 1 0 7270 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_39
timestamp 1676037725
transform 1 0 6646 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_40
timestamp 1676037725
transform 1 0 8272 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_41
timestamp 1676037725
transform 1 0 8736 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_42
timestamp 1676037725
transform 1 0 8140 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_43
timestamp 1676037725
transform 1 0 7676 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_44
timestamp 1676037725
transform 1 0 7024 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_45
timestamp 1676037725
transform 1 0 7488 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_46
timestamp 1676037725
transform 1 0 6892 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_47
timestamp 1676037725
transform 1 0 6428 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_48
timestamp 1676037725
transform 1 0 14512 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_49
timestamp 1676037725
transform 1 0 14976 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_50
timestamp 1676037725
transform 1 0 14380 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_51
timestamp 1676037725
transform 1 0 13916 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_52
timestamp 1676037725
transform 1 0 13264 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_53
timestamp 1676037725
transform 1 0 13728 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_54
timestamp 1676037725
transform 1 0 13132 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_55
timestamp 1676037725
transform 1 0 12668 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_56
timestamp 1676037725
transform 1 0 12016 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_57
timestamp 1676037725
transform 1 0 12480 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_58
timestamp 1676037725
transform 1 0 11884 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_59
timestamp 1676037725
transform 1 0 11420 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_60
timestamp 1676037725
transform 1 0 16006 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_61
timestamp 1676037725
transform 1 0 15382 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_62
timestamp 1676037725
transform 1 0 14758 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_63
timestamp 1676037725
transform 1 0 14134 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_64
timestamp 1676037725
transform 1 0 13510 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_65
timestamp 1676037725
transform 1 0 12886 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_66
timestamp 1676037725
transform 1 0 12262 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_67
timestamp 1676037725
transform 1 0 11638 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_68
timestamp 1676037725
transform 1 0 15760 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_69
timestamp 1676037725
transform 1 0 16224 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_70
timestamp 1676037725
transform 1 0 15628 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_71
timestamp 1676037725
transform 1 0 15164 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_72
timestamp 1676037725
transform 1 0 20998 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_73
timestamp 1676037725
transform 1 0 20374 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_74
timestamp 1676037725
transform 1 0 19750 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_75
timestamp 1676037725
transform 1 0 19126 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_76
timestamp 1676037725
transform 1 0 18502 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_77
timestamp 1676037725
transform 1 0 17878 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_78
timestamp 1676037725
transform 1 0 17254 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_79
timestamp 1676037725
transform 1 0 16630 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_80
timestamp 1676037725
transform 1 0 20752 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_81
timestamp 1676037725
transform 1 0 21216 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_82
timestamp 1676037725
transform 1 0 20620 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_83
timestamp 1676037725
transform 1 0 20156 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_84
timestamp 1676037725
transform 1 0 19504 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_85
timestamp 1676037725
transform 1 0 19968 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_86
timestamp 1676037725
transform 1 0 19372 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_87
timestamp 1676037725
transform 1 0 18908 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_88
timestamp 1676037725
transform 1 0 18256 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_89
timestamp 1676037725
transform 1 0 18720 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_90
timestamp 1676037725
transform 1 0 18124 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_91
timestamp 1676037725
transform 1 0 17660 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_92
timestamp 1676037725
transform 1 0 17008 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_93
timestamp 1676037725
transform 1 0 17472 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_94
timestamp 1676037725
transform 1 0 16876 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_95
timestamp 1676037725
transform 1 0 16412 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_96
timestamp 1676037725
transform 1 0 23494 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_97
timestamp 1676037725
transform 1 0 22870 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_98
timestamp 1676037725
transform 1 0 22246 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_99
timestamp 1676037725
transform 1 0 21622 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_100
timestamp 1676037725
transform 1 0 24496 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_101
timestamp 1676037725
transform 1 0 24960 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_102
timestamp 1676037725
transform 1 0 24364 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_103
timestamp 1676037725
transform 1 0 23900 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_104
timestamp 1676037725
transform 1 0 23248 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_105
timestamp 1676037725
transform 1 0 23712 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_106
timestamp 1676037725
transform 1 0 23116 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_107
timestamp 1676037725
transform 1 0 22652 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_108
timestamp 1676037725
transform 1 0 22000 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_109
timestamp 1676037725
transform 1 0 22464 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_110
timestamp 1676037725
transform 1 0 21868 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_111
timestamp 1676037725
transform 1 0 21404 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_112
timestamp 1676037725
transform 1 0 25990 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_113
timestamp 1676037725
transform 1 0 25366 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_114
timestamp 1676037725
transform 1 0 24742 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_115
timestamp 1676037725
transform 1 0 24118 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_116
timestamp 1676037725
transform 1 0 25744 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_117
timestamp 1676037725
transform 1 0 26208 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_118
timestamp 1676037725
transform 1 0 25612 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_119
timestamp 1676037725
transform 1 0 25148 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_120
timestamp 1676037725
transform 1 0 30736 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_121
timestamp 1676037725
transform 1 0 31200 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_122
timestamp 1676037725
transform 1 0 30604 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_123
timestamp 1676037725
transform 1 0 30140 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_124
timestamp 1676037725
transform 1 0 29488 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_125
timestamp 1676037725
transform 1 0 29952 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_126
timestamp 1676037725
transform 1 0 29356 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_127
timestamp 1676037725
transform 1 0 28892 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_128
timestamp 1676037725
transform 1 0 28240 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_129
timestamp 1676037725
transform 1 0 28704 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_130
timestamp 1676037725
transform 1 0 28108 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_131
timestamp 1676037725
transform 1 0 27644 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_132
timestamp 1676037725
transform 1 0 26992 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_133
timestamp 1676037725
transform 1 0 27456 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_134
timestamp 1676037725
transform 1 0 26860 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_135
timestamp 1676037725
transform 1 0 26396 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_136
timestamp 1676037725
transform 1 0 30982 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_137
timestamp 1676037725
transform 1 0 30358 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_138
timestamp 1676037725
transform 1 0 29734 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_139
timestamp 1676037725
transform 1 0 29110 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_140
timestamp 1676037725
transform 1 0 28486 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_141
timestamp 1676037725
transform 1 0 27862 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_142
timestamp 1676037725
transform 1 0 27238 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_143
timestamp 1676037725
transform 1 0 26614 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_144
timestamp 1676037725
transform 1 0 32230 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_145
timestamp 1676037725
transform 1 0 31606 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_146
timestamp 1676037725
transform 1 0 35728 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_147
timestamp 1676037725
transform 1 0 36192 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_148
timestamp 1676037725
transform 1 0 35596 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_149
timestamp 1676037725
transform 1 0 35132 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_150
timestamp 1676037725
transform 1 0 34480 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_151
timestamp 1676037725
transform 1 0 34944 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_152
timestamp 1676037725
transform 1 0 34348 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_153
timestamp 1676037725
transform 1 0 33884 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_154
timestamp 1676037725
transform 1 0 33232 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_155
timestamp 1676037725
transform 1 0 33696 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_156
timestamp 1676037725
transform 1 0 33100 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_157
timestamp 1676037725
transform 1 0 32636 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_158
timestamp 1676037725
transform 1 0 31984 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_159
timestamp 1676037725
transform 1 0 32448 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_160
timestamp 1676037725
transform 1 0 31852 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_161
timestamp 1676037725
transform 1 0 31388 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_162
timestamp 1676037725
transform 1 0 35974 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_163
timestamp 1676037725
transform 1 0 35350 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_164
timestamp 1676037725
transform 1 0 34726 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_165
timestamp 1676037725
transform 1 0 34102 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_166
timestamp 1676037725
transform 1 0 33478 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_167
timestamp 1676037725
transform 1 0 32854 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_168
timestamp 1676037725
transform 1 0 40966 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_169
timestamp 1676037725
transform 1 0 40342 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_170
timestamp 1676037725
transform 1 0 39718 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_171
timestamp 1676037725
transform 1 0 39094 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_172
timestamp 1676037725
transform 1 0 38470 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_173
timestamp 1676037725
transform 1 0 37846 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_174
timestamp 1676037725
transform 1 0 37222 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_175
timestamp 1676037725
transform 1 0 36598 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_176
timestamp 1676037725
transform 1 0 40720 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_177
timestamp 1676037725
transform 1 0 41184 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_178
timestamp 1676037725
transform 1 0 40588 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_179
timestamp 1676037725
transform 1 0 40124 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_180
timestamp 1676037725
transform 1 0 39472 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_181
timestamp 1676037725
transform 1 0 39936 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_182
timestamp 1676037725
transform 1 0 39340 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_183
timestamp 1676037725
transform 1 0 38876 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_184
timestamp 1676037725
transform 1 0 38224 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_185
timestamp 1676037725
transform 1 0 38688 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_186
timestamp 1676037725
transform 1 0 38092 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_187
timestamp 1676037725
transform 1 0 37628 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_188
timestamp 1676037725
transform 1 0 36976 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_189
timestamp 1676037725
transform 1 0 37440 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_190
timestamp 1676037725
transform 1 0 36844 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_191
timestamp 1676037725
transform 1 0 36380 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_192
timestamp 1676037725
transform 1 0 43216 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_193
timestamp 1676037725
transform 1 0 43680 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_194
timestamp 1676037725
transform 1 0 43084 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_195
timestamp 1676037725
transform 1 0 42620 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_196
timestamp 1676037725
transform 1 0 41968 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_197
timestamp 1676037725
transform 1 0 42432 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_198
timestamp 1676037725
transform 1 0 41836 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_199
timestamp 1676037725
transform 1 0 41372 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_200
timestamp 1676037725
transform 1 0 45712 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_201
timestamp 1676037725
transform 1 0 46176 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_202
timestamp 1676037725
transform 1 0 45580 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_203
timestamp 1676037725
transform 1 0 45116 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_204
timestamp 1676037725
transform 1 0 45958 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_205
timestamp 1676037725
transform 1 0 45334 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_206
timestamp 1676037725
transform 1 0 44710 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_207
timestamp 1676037725
transform 1 0 44086 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_208
timestamp 1676037725
transform 1 0 43462 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_209
timestamp 1676037725
transform 1 0 42838 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_210
timestamp 1676037725
transform 1 0 42214 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_211
timestamp 1676037725
transform 1 0 41590 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_212
timestamp 1676037725
transform 1 0 44464 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_213
timestamp 1676037725
transform 1 0 44928 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_214
timestamp 1676037725
transform 1 0 44332 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_215
timestamp 1676037725
transform 1 0 43868 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_216
timestamp 1676037725
transform 1 0 50950 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_217
timestamp 1676037725
transform 1 0 50326 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_218
timestamp 1676037725
transform 1 0 49702 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_219
timestamp 1676037725
transform 1 0 49078 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_220
timestamp 1676037725
transform 1 0 48454 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_221
timestamp 1676037725
transform 1 0 47830 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_222
timestamp 1676037725
transform 1 0 47206 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_223
timestamp 1676037725
transform 1 0 46582 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_224
timestamp 1676037725
transform 1 0 48208 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_225
timestamp 1676037725
transform 1 0 48672 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_226
timestamp 1676037725
transform 1 0 48076 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_227
timestamp 1676037725
transform 1 0 47612 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_228
timestamp 1676037725
transform 1 0 46960 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_229
timestamp 1676037725
transform 1 0 47424 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_230
timestamp 1676037725
transform 1 0 46828 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_231
timestamp 1676037725
transform 1 0 46364 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_232
timestamp 1676037725
transform 1 0 50704 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_233
timestamp 1676037725
transform 1 0 51168 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_234
timestamp 1676037725
transform 1 0 50572 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_235
timestamp 1676037725
transform 1 0 50108 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_236
timestamp 1676037725
transform 1 0 49456 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_237
timestamp 1676037725
transform 1 0 49920 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_238
timestamp 1676037725
transform 1 0 49324 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_239
timestamp 1676037725
transform 1 0 48860 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_240
timestamp 1676037725
transform 1 0 52198 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_241
timestamp 1676037725
transform 1 0 51574 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_242
timestamp 1676037725
transform 1 0 55696 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_243
timestamp 1676037725
transform 1 0 56160 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_244
timestamp 1676037725
transform 1 0 55564 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_245
timestamp 1676037725
transform 1 0 55100 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_246
timestamp 1676037725
transform 1 0 54448 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_247
timestamp 1676037725
transform 1 0 54912 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_248
timestamp 1676037725
transform 1 0 54316 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_249
timestamp 1676037725
transform 1 0 53852 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_250
timestamp 1676037725
transform 1 0 53200 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_251
timestamp 1676037725
transform 1 0 53664 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_252
timestamp 1676037725
transform 1 0 53068 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_253
timestamp 1676037725
transform 1 0 52604 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_254
timestamp 1676037725
transform 1 0 51952 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_255
timestamp 1676037725
transform 1 0 52416 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_256
timestamp 1676037725
transform 1 0 51820 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_257
timestamp 1676037725
transform 1 0 51356 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_258
timestamp 1676037725
transform 1 0 55942 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_259
timestamp 1676037725
transform 1 0 55318 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_260
timestamp 1676037725
transform 1 0 54694 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_261
timestamp 1676037725
transform 1 0 54070 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_262
timestamp 1676037725
transform 1 0 53446 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_263
timestamp 1676037725
transform 1 0 52822 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_264
timestamp 1676037725
transform 1 0 60934 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_265
timestamp 1676037725
transform 1 0 60310 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_266
timestamp 1676037725
transform 1 0 59686 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_267
timestamp 1676037725
transform 1 0 59062 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_268
timestamp 1676037725
transform 1 0 58438 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_269
timestamp 1676037725
transform 1 0 57814 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_270
timestamp 1676037725
transform 1 0 57190 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_271
timestamp 1676037725
transform 1 0 56566 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_272
timestamp 1676037725
transform 1 0 60688 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_273
timestamp 1676037725
transform 1 0 61152 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_274
timestamp 1676037725
transform 1 0 60556 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_275
timestamp 1676037725
transform 1 0 60092 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_276
timestamp 1676037725
transform 1 0 59440 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_277
timestamp 1676037725
transform 1 0 59904 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_278
timestamp 1676037725
transform 1 0 59308 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_279
timestamp 1676037725
transform 1 0 58844 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_280
timestamp 1676037725
transform 1 0 58192 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_281
timestamp 1676037725
transform 1 0 58656 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_282
timestamp 1676037725
transform 1 0 58060 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_283
timestamp 1676037725
transform 1 0 57596 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_284
timestamp 1676037725
transform 1 0 56944 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_285
timestamp 1676037725
transform 1 0 57408 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_286
timestamp 1676037725
transform 1 0 56812 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_287
timestamp 1676037725
transform 1 0 56348 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_288
timestamp 1676037725
transform 1 0 65926 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_289
timestamp 1676037725
transform 1 0 65302 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_290
timestamp 1676037725
transform 1 0 64678 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_291
timestamp 1676037725
transform 1 0 64054 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_292
timestamp 1676037725
transform 1 0 63430 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_293
timestamp 1676037725
transform 1 0 62806 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_294
timestamp 1676037725
transform 1 0 62182 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_295
timestamp 1676037725
transform 1 0 61558 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_296
timestamp 1676037725
transform 1 0 64432 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_297
timestamp 1676037725
transform 1 0 64896 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_298
timestamp 1676037725
transform 1 0 64300 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_299
timestamp 1676037725
transform 1 0 63836 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_300
timestamp 1676037725
transform 1 0 63184 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_301
timestamp 1676037725
transform 1 0 63648 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_302
timestamp 1676037725
transform 1 0 63052 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_303
timestamp 1676037725
transform 1 0 62588 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_304
timestamp 1676037725
transform 1 0 61936 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_305
timestamp 1676037725
transform 1 0 62400 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_306
timestamp 1676037725
transform 1 0 61804 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_307
timestamp 1676037725
transform 1 0 61340 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_308
timestamp 1676037725
transform 1 0 65680 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_309
timestamp 1676037725
transform 1 0 66144 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_310
timestamp 1676037725
transform 1 0 65548 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_311
timestamp 1676037725
transform 1 0 65084 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_312
timestamp 1676037725
transform 1 0 70918 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_313
timestamp 1676037725
transform 1 0 70294 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_314
timestamp 1676037725
transform 1 0 69670 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_315
timestamp 1676037725
transform 1 0 69046 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_316
timestamp 1676037725
transform 1 0 70672 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_317
timestamp 1676037725
transform 1 0 71136 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_318
timestamp 1676037725
transform 1 0 70540 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_319
timestamp 1676037725
transform 1 0 70076 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_320
timestamp 1676037725
transform 1 0 69424 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_321
timestamp 1676037725
transform 1 0 69888 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_322
timestamp 1676037725
transform 1 0 69292 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_323
timestamp 1676037725
transform 1 0 68828 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_324
timestamp 1676037725
transform 1 0 68176 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_325
timestamp 1676037725
transform 1 0 68640 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_326
timestamp 1676037725
transform 1 0 68044 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_327
timestamp 1676037725
transform 1 0 67580 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_328
timestamp 1676037725
transform 1 0 66928 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_329
timestamp 1676037725
transform 1 0 67392 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_330
timestamp 1676037725
transform 1 0 66796 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_331
timestamp 1676037725
transform 1 0 66332 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_332
timestamp 1676037725
transform 1 0 68422 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_333
timestamp 1676037725
transform 1 0 67798 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_334
timestamp 1676037725
transform 1 0 67174 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_335
timestamp 1676037725
transform 1 0 66550 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_336
timestamp 1676037725
transform 1 0 73414 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_337
timestamp 1676037725
transform 1 0 72790 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_338
timestamp 1676037725
transform 1 0 72166 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_339
timestamp 1676037725
transform 1 0 71542 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_340
timestamp 1676037725
transform 1 0 75910 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_341
timestamp 1676037725
transform 1 0 75286 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_342
timestamp 1676037725
transform 1 0 75664 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_343
timestamp 1676037725
transform 1 0 76128 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_344
timestamp 1676037725
transform 1 0 75532 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_345
timestamp 1676037725
transform 1 0 75068 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_346
timestamp 1676037725
transform 1 0 74416 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_347
timestamp 1676037725
transform 1 0 74880 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_348
timestamp 1676037725
transform 1 0 74284 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_349
timestamp 1676037725
transform 1 0 73820 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_350
timestamp 1676037725
transform 1 0 73168 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_351
timestamp 1676037725
transform 1 0 73632 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_352
timestamp 1676037725
transform 1 0 73036 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_353
timestamp 1676037725
transform 1 0 72572 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_354
timestamp 1676037725
transform 1 0 71920 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_355
timestamp 1676037725
transform 1 0 72384 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_356
timestamp 1676037725
transform 1 0 71788 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_357
timestamp 1676037725
transform 1 0 71324 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_358
timestamp 1676037725
transform 1 0 74662 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_359
timestamp 1676037725
transform 1 0 74038 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_360
timestamp 1676037725
transform 1 0 80656 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_361
timestamp 1676037725
transform 1 0 81120 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_362
timestamp 1676037725
transform 1 0 80524 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_363
timestamp 1676037725
transform 1 0 80060 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_364
timestamp 1676037725
transform 1 0 79408 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_365
timestamp 1676037725
transform 1 0 79872 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_366
timestamp 1676037725
transform 1 0 79276 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_367
timestamp 1676037725
transform 1 0 78812 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_368
timestamp 1676037725
transform 1 0 78160 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_369
timestamp 1676037725
transform 1 0 78624 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_370
timestamp 1676037725
transform 1 0 78028 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_371
timestamp 1676037725
transform 1 0 77564 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_372
timestamp 1676037725
transform 1 0 76912 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_373
timestamp 1676037725
transform 1 0 77376 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_374
timestamp 1676037725
transform 1 0 76780 0 1 92
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_375
timestamp 1676037725
transform 1 0 76316 0 1 216
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_376
timestamp 1676037725
transform 1 0 80902 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_377
timestamp 1676037725
transform 1 0 80278 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_378
timestamp 1676037725
transform 1 0 79654 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_379
timestamp 1676037725
transform 1 0 79030 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_380
timestamp 1676037725
transform 1 0 78406 0 1 742
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_381
timestamp 1676037725
transform 1 0 77782 0 1 618
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_382
timestamp 1676037725
transform 1 0 77158 0 1 494
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_26  sky130_sram_2kbyte_1rw1r_32x512_8_contact_26_383
timestamp 1676037725
transform 1 0 76534 0 1 370
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_0
timestamp 1676037725
transform 1 0 5775 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_1
timestamp 1676037725
transform 1 0 6239 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_2
timestamp 1676037725
transform 1 0 5643 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_3
timestamp 1676037725
transform 1 0 5179 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_4
timestamp 1676037725
transform 1 0 4527 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_5
timestamp 1676037725
transform 1 0 4991 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_6
timestamp 1676037725
transform 1 0 4395 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_7
timestamp 1676037725
transform 1 0 3931 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_8
timestamp 1676037725
transform 1 0 3279 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_9
timestamp 1676037725
transform 1 0 3743 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_10
timestamp 1676037725
transform 1 0 3147 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_11
timestamp 1676037725
transform 1 0 2683 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_12
timestamp 1676037725
transform 1 0 2031 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_13
timestamp 1676037725
transform 1 0 2495 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_14
timestamp 1676037725
transform 1 0 1899 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_15
timestamp 1676037725
transform 1 0 1435 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_16
timestamp 1676037725
transform 1 0 4773 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_17
timestamp 1676037725
transform 1 0 4149 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_18
timestamp 1676037725
transform 1 0 3525 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_19
timestamp 1676037725
transform 1 0 2901 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_20
timestamp 1676037725
transform 1 0 2277 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_21
timestamp 1676037725
transform 1 0 1653 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_22
timestamp 1676037725
transform 1 0 6021 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_23
timestamp 1676037725
transform 1 0 5397 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_24
timestamp 1676037725
transform 1 0 10767 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_25
timestamp 1676037725
transform 1 0 11231 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_26
timestamp 1676037725
transform 1 0 10635 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_27
timestamp 1676037725
transform 1 0 10171 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_28
timestamp 1676037725
transform 1 0 9519 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_29
timestamp 1676037725
transform 1 0 9983 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_30
timestamp 1676037725
transform 1 0 9387 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_31
timestamp 1676037725
transform 1 0 8923 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_32
timestamp 1676037725
transform 1 0 11013 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_33
timestamp 1676037725
transform 1 0 10389 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_34
timestamp 1676037725
transform 1 0 9765 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_35
timestamp 1676037725
transform 1 0 9141 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_36
timestamp 1676037725
transform 1 0 8517 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_37
timestamp 1676037725
transform 1 0 7893 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_38
timestamp 1676037725
transform 1 0 7269 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_39
timestamp 1676037725
transform 1 0 6645 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_40
timestamp 1676037725
transform 1 0 8271 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_41
timestamp 1676037725
transform 1 0 8735 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_42
timestamp 1676037725
transform 1 0 8139 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_43
timestamp 1676037725
transform 1 0 7675 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_44
timestamp 1676037725
transform 1 0 7023 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_45
timestamp 1676037725
transform 1 0 7487 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_46
timestamp 1676037725
transform 1 0 6891 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_47
timestamp 1676037725
transform 1 0 6427 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_48
timestamp 1676037725
transform 1 0 14511 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_49
timestamp 1676037725
transform 1 0 14975 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_50
timestamp 1676037725
transform 1 0 14379 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_51
timestamp 1676037725
transform 1 0 13915 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_52
timestamp 1676037725
transform 1 0 13263 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_53
timestamp 1676037725
transform 1 0 13727 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_54
timestamp 1676037725
transform 1 0 13131 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_55
timestamp 1676037725
transform 1 0 12667 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_56
timestamp 1676037725
transform 1 0 12015 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_57
timestamp 1676037725
transform 1 0 12479 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_58
timestamp 1676037725
transform 1 0 11883 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_59
timestamp 1676037725
transform 1 0 11419 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_60
timestamp 1676037725
transform 1 0 16005 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_61
timestamp 1676037725
transform 1 0 15381 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_62
timestamp 1676037725
transform 1 0 14757 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_63
timestamp 1676037725
transform 1 0 14133 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_64
timestamp 1676037725
transform 1 0 13509 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_65
timestamp 1676037725
transform 1 0 12885 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_66
timestamp 1676037725
transform 1 0 12261 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_67
timestamp 1676037725
transform 1 0 11637 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_68
timestamp 1676037725
transform 1 0 15759 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_69
timestamp 1676037725
transform 1 0 16223 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_70
timestamp 1676037725
transform 1 0 15627 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_71
timestamp 1676037725
transform 1 0 15163 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_72
timestamp 1676037725
transform 1 0 20997 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_73
timestamp 1676037725
transform 1 0 20373 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_74
timestamp 1676037725
transform 1 0 19749 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_75
timestamp 1676037725
transform 1 0 19125 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_76
timestamp 1676037725
transform 1 0 18501 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_77
timestamp 1676037725
transform 1 0 17877 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_78
timestamp 1676037725
transform 1 0 17253 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_79
timestamp 1676037725
transform 1 0 16629 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_80
timestamp 1676037725
transform 1 0 20751 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_81
timestamp 1676037725
transform 1 0 21215 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_82
timestamp 1676037725
transform 1 0 20619 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_83
timestamp 1676037725
transform 1 0 20155 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_84
timestamp 1676037725
transform 1 0 19503 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_85
timestamp 1676037725
transform 1 0 19967 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_86
timestamp 1676037725
transform 1 0 19371 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_87
timestamp 1676037725
transform 1 0 18907 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_88
timestamp 1676037725
transform 1 0 18255 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_89
timestamp 1676037725
transform 1 0 18719 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_90
timestamp 1676037725
transform 1 0 18123 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_91
timestamp 1676037725
transform 1 0 17659 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_92
timestamp 1676037725
transform 1 0 17007 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_93
timestamp 1676037725
transform 1 0 17471 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_94
timestamp 1676037725
transform 1 0 16875 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_95
timestamp 1676037725
transform 1 0 16411 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_96
timestamp 1676037725
transform 1 0 23493 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_97
timestamp 1676037725
transform 1 0 22869 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_98
timestamp 1676037725
transform 1 0 22245 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_99
timestamp 1676037725
transform 1 0 21621 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_100
timestamp 1676037725
transform 1 0 24495 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_101
timestamp 1676037725
transform 1 0 24959 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_102
timestamp 1676037725
transform 1 0 24363 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_103
timestamp 1676037725
transform 1 0 23899 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_104
timestamp 1676037725
transform 1 0 23247 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_105
timestamp 1676037725
transform 1 0 23711 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_106
timestamp 1676037725
transform 1 0 23115 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_107
timestamp 1676037725
transform 1 0 22651 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_108
timestamp 1676037725
transform 1 0 21999 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_109
timestamp 1676037725
transform 1 0 22463 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_110
timestamp 1676037725
transform 1 0 21867 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_111
timestamp 1676037725
transform 1 0 21403 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_112
timestamp 1676037725
transform 1 0 25989 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_113
timestamp 1676037725
transform 1 0 25365 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_114
timestamp 1676037725
transform 1 0 24741 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_115
timestamp 1676037725
transform 1 0 24117 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_116
timestamp 1676037725
transform 1 0 25743 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_117
timestamp 1676037725
transform 1 0 26207 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_118
timestamp 1676037725
transform 1 0 25611 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_119
timestamp 1676037725
transform 1 0 25147 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_120
timestamp 1676037725
transform 1 0 30735 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_121
timestamp 1676037725
transform 1 0 31199 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_122
timestamp 1676037725
transform 1 0 30603 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_123
timestamp 1676037725
transform 1 0 30139 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_124
timestamp 1676037725
transform 1 0 29487 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_125
timestamp 1676037725
transform 1 0 29951 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_126
timestamp 1676037725
transform 1 0 29355 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_127
timestamp 1676037725
transform 1 0 28891 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_128
timestamp 1676037725
transform 1 0 28239 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_129
timestamp 1676037725
transform 1 0 28703 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_130
timestamp 1676037725
transform 1 0 28107 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_131
timestamp 1676037725
transform 1 0 27643 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_132
timestamp 1676037725
transform 1 0 26991 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_133
timestamp 1676037725
transform 1 0 27455 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_134
timestamp 1676037725
transform 1 0 26859 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_135
timestamp 1676037725
transform 1 0 26395 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_136
timestamp 1676037725
transform 1 0 30981 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_137
timestamp 1676037725
transform 1 0 30357 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_138
timestamp 1676037725
transform 1 0 29733 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_139
timestamp 1676037725
transform 1 0 29109 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_140
timestamp 1676037725
transform 1 0 28485 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_141
timestamp 1676037725
transform 1 0 27861 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_142
timestamp 1676037725
transform 1 0 27237 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_143
timestamp 1676037725
transform 1 0 26613 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_144
timestamp 1676037725
transform 1 0 32229 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_145
timestamp 1676037725
transform 1 0 31605 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_146
timestamp 1676037725
transform 1 0 35727 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_147
timestamp 1676037725
transform 1 0 36191 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_148
timestamp 1676037725
transform 1 0 35595 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_149
timestamp 1676037725
transform 1 0 35131 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_150
timestamp 1676037725
transform 1 0 34479 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_151
timestamp 1676037725
transform 1 0 34943 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_152
timestamp 1676037725
transform 1 0 34347 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_153
timestamp 1676037725
transform 1 0 33883 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_154
timestamp 1676037725
transform 1 0 33231 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_155
timestamp 1676037725
transform 1 0 33695 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_156
timestamp 1676037725
transform 1 0 33099 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_157
timestamp 1676037725
transform 1 0 32635 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_158
timestamp 1676037725
transform 1 0 31983 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_159
timestamp 1676037725
transform 1 0 32447 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_160
timestamp 1676037725
transform 1 0 31851 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_161
timestamp 1676037725
transform 1 0 31387 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_162
timestamp 1676037725
transform 1 0 35973 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_163
timestamp 1676037725
transform 1 0 35349 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_164
timestamp 1676037725
transform 1 0 34725 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_165
timestamp 1676037725
transform 1 0 34101 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_166
timestamp 1676037725
transform 1 0 33477 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_167
timestamp 1676037725
transform 1 0 32853 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_168
timestamp 1676037725
transform 1 0 40965 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_169
timestamp 1676037725
transform 1 0 40341 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_170
timestamp 1676037725
transform 1 0 39717 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_171
timestamp 1676037725
transform 1 0 39093 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_172
timestamp 1676037725
transform 1 0 38469 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_173
timestamp 1676037725
transform 1 0 37845 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_174
timestamp 1676037725
transform 1 0 37221 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_175
timestamp 1676037725
transform 1 0 36597 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_176
timestamp 1676037725
transform 1 0 40719 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_177
timestamp 1676037725
transform 1 0 41183 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_178
timestamp 1676037725
transform 1 0 40587 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_179
timestamp 1676037725
transform 1 0 40123 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_180
timestamp 1676037725
transform 1 0 39471 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_181
timestamp 1676037725
transform 1 0 39935 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_182
timestamp 1676037725
transform 1 0 39339 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_183
timestamp 1676037725
transform 1 0 38875 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_184
timestamp 1676037725
transform 1 0 38223 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_185
timestamp 1676037725
transform 1 0 38687 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_186
timestamp 1676037725
transform 1 0 38091 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_187
timestamp 1676037725
transform 1 0 37627 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_188
timestamp 1676037725
transform 1 0 36975 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_189
timestamp 1676037725
transform 1 0 37439 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_190
timestamp 1676037725
transform 1 0 36843 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_191
timestamp 1676037725
transform 1 0 36379 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_192
timestamp 1676037725
transform 1 0 43215 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_193
timestamp 1676037725
transform 1 0 43679 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_194
timestamp 1676037725
transform 1 0 43083 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_195
timestamp 1676037725
transform 1 0 42619 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_196
timestamp 1676037725
transform 1 0 41967 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_197
timestamp 1676037725
transform 1 0 42431 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_198
timestamp 1676037725
transform 1 0 41835 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_199
timestamp 1676037725
transform 1 0 41371 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_200
timestamp 1676037725
transform 1 0 45711 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_201
timestamp 1676037725
transform 1 0 46175 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_202
timestamp 1676037725
transform 1 0 45579 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_203
timestamp 1676037725
transform 1 0 45115 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_204
timestamp 1676037725
transform 1 0 45957 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_205
timestamp 1676037725
transform 1 0 45333 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_206
timestamp 1676037725
transform 1 0 44709 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_207
timestamp 1676037725
transform 1 0 44085 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_208
timestamp 1676037725
transform 1 0 43461 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_209
timestamp 1676037725
transform 1 0 42837 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_210
timestamp 1676037725
transform 1 0 42213 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_211
timestamp 1676037725
transform 1 0 41589 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_212
timestamp 1676037725
transform 1 0 44463 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_213
timestamp 1676037725
transform 1 0 44927 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_214
timestamp 1676037725
transform 1 0 44331 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_215
timestamp 1676037725
transform 1 0 43867 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_216
timestamp 1676037725
transform 1 0 50949 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_217
timestamp 1676037725
transform 1 0 50325 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_218
timestamp 1676037725
transform 1 0 49701 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_219
timestamp 1676037725
transform 1 0 49077 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_220
timestamp 1676037725
transform 1 0 48453 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_221
timestamp 1676037725
transform 1 0 47829 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_222
timestamp 1676037725
transform 1 0 47205 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_223
timestamp 1676037725
transform 1 0 46581 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_224
timestamp 1676037725
transform 1 0 48207 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_225
timestamp 1676037725
transform 1 0 48671 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_226
timestamp 1676037725
transform 1 0 48075 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_227
timestamp 1676037725
transform 1 0 47611 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_228
timestamp 1676037725
transform 1 0 46959 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_229
timestamp 1676037725
transform 1 0 47423 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_230
timestamp 1676037725
transform 1 0 46827 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_231
timestamp 1676037725
transform 1 0 46363 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_232
timestamp 1676037725
transform 1 0 50703 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_233
timestamp 1676037725
transform 1 0 51167 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_234
timestamp 1676037725
transform 1 0 50571 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_235
timestamp 1676037725
transform 1 0 50107 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_236
timestamp 1676037725
transform 1 0 49455 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_237
timestamp 1676037725
transform 1 0 49919 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_238
timestamp 1676037725
transform 1 0 49323 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_239
timestamp 1676037725
transform 1 0 48859 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_240
timestamp 1676037725
transform 1 0 52197 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_241
timestamp 1676037725
transform 1 0 51573 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_242
timestamp 1676037725
transform 1 0 55695 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_243
timestamp 1676037725
transform 1 0 56159 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_244
timestamp 1676037725
transform 1 0 55563 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_245
timestamp 1676037725
transform 1 0 55099 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_246
timestamp 1676037725
transform 1 0 54447 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_247
timestamp 1676037725
transform 1 0 54911 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_248
timestamp 1676037725
transform 1 0 54315 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_249
timestamp 1676037725
transform 1 0 53851 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_250
timestamp 1676037725
transform 1 0 53199 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_251
timestamp 1676037725
transform 1 0 53663 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_252
timestamp 1676037725
transform 1 0 53067 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_253
timestamp 1676037725
transform 1 0 52603 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_254
timestamp 1676037725
transform 1 0 51951 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_255
timestamp 1676037725
transform 1 0 52415 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_256
timestamp 1676037725
transform 1 0 51819 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_257
timestamp 1676037725
transform 1 0 51355 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_258
timestamp 1676037725
transform 1 0 55941 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_259
timestamp 1676037725
transform 1 0 55317 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_260
timestamp 1676037725
transform 1 0 54693 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_261
timestamp 1676037725
transform 1 0 54069 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_262
timestamp 1676037725
transform 1 0 53445 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_263
timestamp 1676037725
transform 1 0 52821 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_264
timestamp 1676037725
transform 1 0 60933 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_265
timestamp 1676037725
transform 1 0 60309 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_266
timestamp 1676037725
transform 1 0 59685 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_267
timestamp 1676037725
transform 1 0 59061 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_268
timestamp 1676037725
transform 1 0 58437 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_269
timestamp 1676037725
transform 1 0 57813 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_270
timestamp 1676037725
transform 1 0 57189 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_271
timestamp 1676037725
transform 1 0 56565 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_272
timestamp 1676037725
transform 1 0 60687 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_273
timestamp 1676037725
transform 1 0 61151 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_274
timestamp 1676037725
transform 1 0 60555 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_275
timestamp 1676037725
transform 1 0 60091 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_276
timestamp 1676037725
transform 1 0 59439 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_277
timestamp 1676037725
transform 1 0 59903 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_278
timestamp 1676037725
transform 1 0 59307 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_279
timestamp 1676037725
transform 1 0 58843 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_280
timestamp 1676037725
transform 1 0 58191 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_281
timestamp 1676037725
transform 1 0 58655 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_282
timestamp 1676037725
transform 1 0 58059 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_283
timestamp 1676037725
transform 1 0 57595 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_284
timestamp 1676037725
transform 1 0 56943 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_285
timestamp 1676037725
transform 1 0 57407 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_286
timestamp 1676037725
transform 1 0 56811 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_287
timestamp 1676037725
transform 1 0 56347 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_288
timestamp 1676037725
transform 1 0 65925 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_289
timestamp 1676037725
transform 1 0 65301 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_290
timestamp 1676037725
transform 1 0 64677 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_291
timestamp 1676037725
transform 1 0 64053 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_292
timestamp 1676037725
transform 1 0 63429 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_293
timestamp 1676037725
transform 1 0 62805 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_294
timestamp 1676037725
transform 1 0 62181 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_295
timestamp 1676037725
transform 1 0 61557 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_296
timestamp 1676037725
transform 1 0 64431 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_297
timestamp 1676037725
transform 1 0 64895 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_298
timestamp 1676037725
transform 1 0 64299 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_299
timestamp 1676037725
transform 1 0 63835 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_300
timestamp 1676037725
transform 1 0 63183 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_301
timestamp 1676037725
transform 1 0 63647 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_302
timestamp 1676037725
transform 1 0 63051 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_303
timestamp 1676037725
transform 1 0 62587 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_304
timestamp 1676037725
transform 1 0 61935 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_305
timestamp 1676037725
transform 1 0 62399 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_306
timestamp 1676037725
transform 1 0 61803 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_307
timestamp 1676037725
transform 1 0 61339 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_308
timestamp 1676037725
transform 1 0 65679 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_309
timestamp 1676037725
transform 1 0 66143 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_310
timestamp 1676037725
transform 1 0 65547 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_311
timestamp 1676037725
transform 1 0 65083 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_312
timestamp 1676037725
transform 1 0 70917 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_313
timestamp 1676037725
transform 1 0 70293 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_314
timestamp 1676037725
transform 1 0 69669 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_315
timestamp 1676037725
transform 1 0 69045 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_316
timestamp 1676037725
transform 1 0 70671 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_317
timestamp 1676037725
transform 1 0 71135 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_318
timestamp 1676037725
transform 1 0 70539 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_319
timestamp 1676037725
transform 1 0 70075 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_320
timestamp 1676037725
transform 1 0 69423 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_321
timestamp 1676037725
transform 1 0 69887 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_322
timestamp 1676037725
transform 1 0 69291 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_323
timestamp 1676037725
transform 1 0 68827 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_324
timestamp 1676037725
transform 1 0 68175 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_325
timestamp 1676037725
transform 1 0 68639 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_326
timestamp 1676037725
transform 1 0 68043 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_327
timestamp 1676037725
transform 1 0 67579 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_328
timestamp 1676037725
transform 1 0 66927 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_329
timestamp 1676037725
transform 1 0 67391 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_330
timestamp 1676037725
transform 1 0 66795 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_331
timestamp 1676037725
transform 1 0 66331 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_332
timestamp 1676037725
transform 1 0 68421 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_333
timestamp 1676037725
transform 1 0 67797 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_334
timestamp 1676037725
transform 1 0 67173 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_335
timestamp 1676037725
transform 1 0 66549 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_336
timestamp 1676037725
transform 1 0 73413 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_337
timestamp 1676037725
transform 1 0 72789 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_338
timestamp 1676037725
transform 1 0 72165 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_339
timestamp 1676037725
transform 1 0 71541 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_340
timestamp 1676037725
transform 1 0 75909 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_341
timestamp 1676037725
transform 1 0 75285 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_342
timestamp 1676037725
transform 1 0 75663 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_343
timestamp 1676037725
transform 1 0 76127 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_344
timestamp 1676037725
transform 1 0 75531 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_345
timestamp 1676037725
transform 1 0 75067 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_346
timestamp 1676037725
transform 1 0 74415 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_347
timestamp 1676037725
transform 1 0 74879 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_348
timestamp 1676037725
transform 1 0 74283 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_349
timestamp 1676037725
transform 1 0 73819 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_350
timestamp 1676037725
transform 1 0 73167 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_351
timestamp 1676037725
transform 1 0 73631 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_352
timestamp 1676037725
transform 1 0 73035 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_353
timestamp 1676037725
transform 1 0 72571 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_354
timestamp 1676037725
transform 1 0 71919 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_355
timestamp 1676037725
transform 1 0 72383 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_356
timestamp 1676037725
transform 1 0 71787 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_357
timestamp 1676037725
transform 1 0 71323 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_358
timestamp 1676037725
transform 1 0 74661 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_359
timestamp 1676037725
transform 1 0 74037 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_360
timestamp 1676037725
transform 1 0 80655 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_361
timestamp 1676037725
transform 1 0 81119 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_362
timestamp 1676037725
transform 1 0 80523 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_363
timestamp 1676037725
transform 1 0 80059 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_364
timestamp 1676037725
transform 1 0 79407 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_365
timestamp 1676037725
transform 1 0 79871 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_366
timestamp 1676037725
transform 1 0 79275 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_367
timestamp 1676037725
transform 1 0 78811 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_368
timestamp 1676037725
transform 1 0 78159 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_369
timestamp 1676037725
transform 1 0 78623 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_370
timestamp 1676037725
transform 1 0 78027 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_371
timestamp 1676037725
transform 1 0 77563 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_372
timestamp 1676037725
transform 1 0 76911 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_373
timestamp 1676037725
transform 1 0 77375 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_374
timestamp 1676037725
transform 1 0 76779 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_375
timestamp 1676037725
transform 1 0 76315 0 1 211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_376
timestamp 1676037725
transform 1 0 80901 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_377
timestamp 1676037725
transform 1 0 80277 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_378
timestamp 1676037725
transform 1 0 79653 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_379
timestamp 1676037725
transform 1 0 79029 0 1 365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_380
timestamp 1676037725
transform 1 0 78405 0 1 737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_381
timestamp 1676037725
transform 1 0 77781 0 1 613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_382
timestamp 1676037725
transform 1 0 77157 0 1 489
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_27  sky130_sram_2kbyte_1rw1r_32x512_8_contact_27_383
timestamp 1676037725
transform 1 0 76533 0 1 365
box 0 0 1 1
<< labels >>
rlabel metal3 s 0 372 81246 432 4 sel_0
port 1 nsew
rlabel metal3 s 0 496 81246 556 4 sel_1
port 2 nsew
rlabel metal3 s 0 620 81246 680 4 sel_2
port 3 nsew
rlabel metal3 s 0 744 81246 804 4 sel_3
port 4 nsew
rlabel metal3 s 56861 1482 56959 1580 4 gnd
port 5 nsew
rlabel metal3 s 26909 1482 27007 1580 4 gnd
port 5 nsew
rlabel metal3 s 5693 1482 5791 1580 4 gnd
port 5 nsew
rlabel metal3 s 5742 1531 5742 1531 4 gnd
rlabel metal3 s 26958 1531 26958 1531 4 gnd
rlabel metal3 s 60605 1482 60703 1580 4 gnd
port 5 nsew
rlabel metal3 s 60654 1531 60654 1531 4 gnd
rlabel metal3 s 31901 1482 31999 1580 4 gnd
port 5 nsew
rlabel metal3 s 3197 1482 3295 1580 4 gnd
port 5 nsew
rlabel metal3 s 3246 1531 3246 1531 4 gnd
rlabel metal3 s 23165 1482 23263 1580 4 gnd
port 5 nsew
rlabel metal3 s 73085 1482 73183 1580 4 gnd
port 5 nsew
rlabel metal3 s 45629 1482 45727 1580 4 gnd
port 5 nsew
rlabel metal3 s 45678 1531 45678 1531 4 gnd
rlabel metal3 s 74333 1482 74431 1580 4 gnd
port 5 nsew
rlabel metal3 s 64349 1482 64447 1580 4 gnd
port 5 nsew
rlabel metal3 s 53117 1482 53215 1580 4 gnd
port 5 nsew
rlabel metal3 s 41885 1482 41983 1580 4 gnd
port 5 nsew
rlabel metal3 s 41934 1531 41934 1531 4 gnd
rlabel metal3 s 44381 1482 44479 1580 4 gnd
port 5 nsew
rlabel metal3 s 29405 1482 29503 1580 4 gnd
port 5 nsew
rlabel metal3 s 34397 1482 34495 1580 4 gnd
port 5 nsew
rlabel metal3 s 34446 1531 34446 1531 4 gnd
rlabel metal3 s 24413 1482 24511 1580 4 gnd
port 5 nsew
rlabel metal3 s 24462 1531 24462 1531 4 gnd
rlabel metal3 s 39389 1482 39487 1580 4 gnd
port 5 nsew
rlabel metal3 s 20669 1482 20767 1580 4 gnd
port 5 nsew
rlabel metal3 s 20718 1531 20718 1531 4 gnd
rlabel metal3 s 69341 1482 69439 1580 4 gnd
port 5 nsew
rlabel metal3 s 16925 1482 17023 1580 4 gnd
port 5 nsew
rlabel metal3 s 10685 1482 10783 1580 4 gnd
port 5 nsew
rlabel metal3 s 10734 1531 10734 1531 4 gnd
rlabel metal3 s 21917 1482 22015 1580 4 gnd
port 5 nsew
rlabel metal3 s 1949 1482 2047 1580 4 gnd
port 5 nsew
rlabel metal3 s 1998 1531 1998 1531 4 gnd
rlabel metal3 s 48125 1482 48223 1580 4 gnd
port 5 nsew
rlabel metal3 s 50621 1482 50719 1580 4 gnd
port 5 nsew
rlabel metal3 s 70589 1482 70687 1580 4 gnd
port 5 nsew
rlabel metal3 s 63101 1482 63199 1580 4 gnd
port 5 nsew
rlabel metal3 s 6941 1482 7039 1580 4 gnd
port 5 nsew
rlabel metal3 s 66845 1482 66943 1580 4 gnd
port 5 nsew
rlabel metal3 s 8189 1482 8287 1580 4 gnd
port 5 nsew
rlabel metal3 s 59357 1482 59455 1580 4 gnd
port 5 nsew
rlabel metal3 s 79325 1482 79423 1580 4 gnd
port 5 nsew
rlabel metal3 s 75581 1482 75679 1580 4 gnd
port 5 nsew
rlabel metal3 s 75630 1531 75630 1531 4 gnd
rlabel metal3 s 38141 1482 38239 1580 4 gnd
port 5 nsew
rlabel metal3 s 30653 1482 30751 1580 4 gnd
port 5 nsew
rlabel metal3 s 30702 1531 30702 1531 4 gnd
rlabel metal3 s 38190 1531 38190 1531 4 gnd
rlabel metal3 s 33149 1482 33247 1580 4 gnd
port 5 nsew
rlabel metal3 s 40637 1482 40735 1580 4 gnd
port 5 nsew
rlabel metal3 s 65597 1482 65695 1580 4 gnd
port 5 nsew
rlabel metal3 s 80573 1482 80671 1580 4 gnd
port 5 nsew
rlabel metal3 s 28157 1482 28255 1580 4 gnd
port 5 nsew
rlabel metal3 s 68093 1482 68191 1580 4 gnd
port 5 nsew
rlabel metal3 s 68142 1531 68142 1531 4 gnd
rlabel metal3 s 71837 1482 71935 1580 4 gnd
port 5 nsew
rlabel metal3 s 25661 1482 25759 1580 4 gnd
port 5 nsew
rlabel metal3 s 76829 1482 76927 1580 4 gnd
port 5 nsew
rlabel metal3 s 11933 1482 12031 1580 4 gnd
port 5 nsew
rlabel metal3 s 46877 1482 46975 1580 4 gnd
port 5 nsew
rlabel metal3 s 14429 1482 14527 1580 4 gnd
port 5 nsew
rlabel metal3 s 14478 1531 14478 1531 4 gnd
rlabel metal3 s 13181 1482 13279 1580 4 gnd
port 5 nsew
rlabel metal3 s 4445 1482 4543 1580 4 gnd
port 5 nsew
rlabel metal3 s 4494 1531 4494 1531 4 gnd
rlabel metal3 s 18173 1482 18271 1580 4 gnd
port 5 nsew
rlabel metal3 s 18222 1531 18222 1531 4 gnd
rlabel metal3 s 58109 1482 58207 1580 4 gnd
port 5 nsew
rlabel metal3 s 36893 1482 36991 1580 4 gnd
port 5 nsew
rlabel metal3 s 49373 1482 49471 1580 4 gnd
port 5 nsew
rlabel metal3 s 78077 1482 78175 1580 4 gnd
port 5 nsew
rlabel metal3 s 51869 1482 51967 1580 4 gnd
port 5 nsew
rlabel metal3 s 51918 1531 51918 1531 4 gnd
rlabel metal3 s 19421 1482 19519 1580 4 gnd
port 5 nsew
rlabel metal3 s 15677 1482 15775 1580 4 gnd
port 5 nsew
rlabel metal3 s 54365 1482 54463 1580 4 gnd
port 5 nsew
rlabel metal3 s 9437 1482 9535 1580 4 gnd
port 5 nsew
rlabel metal3 s 61853 1482 61951 1580 4 gnd
port 5 nsew
rlabel metal3 s 35645 1482 35743 1580 4 gnd
port 5 nsew
rlabel metal3 s 55613 1482 55711 1580 4 gnd
port 5 nsew
rlabel metal3 s 43133 1482 43231 1580 4 gnd
port 5 nsew
rlabel metal1 s 61358 248 61386 868 4 bl_out_24
port 6 nsew
rlabel metal1 s 63854 248 63882 868 4 bl_out_25
port 7 nsew
rlabel metal1 s 66350 248 66378 868 4 bl_out_26
port 8 nsew
rlabel metal1 s 68846 248 68874 868 4 bl_out_27
port 9 nsew
rlabel metal1 s 71342 248 71370 868 4 bl_out_28
port 10 nsew
rlabel metal1 s 73838 248 73866 868 4 bl_out_29
port 11 nsew
rlabel metal1 s 76334 248 76362 868 4 bl_out_30
port 12 nsew
rlabel metal1 s 78830 248 78858 868 4 bl_out_31
port 13 nsew
rlabel metal1 s 61358 2128 61386 2184 4 bl_96
port 14 nsew
rlabel metal1 s 61822 2128 61850 2184 4 br_96
port 15 nsew
rlabel metal1 s 62418 2128 62446 2184 4 bl_97
port 16 nsew
rlabel metal1 s 61954 2128 61982 2184 4 br_97
port 17 nsew
rlabel metal1 s 62606 2128 62634 2184 4 bl_98
port 18 nsew
rlabel metal1 s 63070 2128 63098 2184 4 br_98
port 19 nsew
rlabel metal1 s 63666 2128 63694 2184 4 bl_99
port 20 nsew
rlabel metal1 s 63202 2128 63230 2184 4 br_99
port 21 nsew
rlabel metal1 s 63854 2128 63882 2184 4 bl_100
port 22 nsew
rlabel metal1 s 64318 2128 64346 2184 4 br_100
port 23 nsew
rlabel metal1 s 64914 2128 64942 2184 4 bl_101
port 24 nsew
rlabel metal1 s 64450 2128 64478 2184 4 br_101
port 25 nsew
rlabel metal1 s 65102 2128 65130 2184 4 bl_102
port 26 nsew
rlabel metal1 s 65566 2128 65594 2184 4 br_102
port 27 nsew
rlabel metal1 s 66162 2128 66190 2184 4 bl_103
port 28 nsew
rlabel metal1 s 65698 2128 65726 2184 4 br_103
port 29 nsew
rlabel metal1 s 66350 2128 66378 2184 4 bl_104
port 30 nsew
rlabel metal1 s 66814 2128 66842 2184 4 br_104
port 31 nsew
rlabel metal1 s 67410 2128 67438 2184 4 bl_105
port 32 nsew
rlabel metal1 s 66946 2128 66974 2184 4 br_105
port 33 nsew
rlabel metal1 s 67598 2128 67626 2184 4 bl_106
port 34 nsew
rlabel metal1 s 68062 2128 68090 2184 4 br_106
port 35 nsew
rlabel metal1 s 68658 2128 68686 2184 4 bl_107
port 36 nsew
rlabel metal1 s 68194 2128 68222 2184 4 br_107
port 37 nsew
rlabel metal1 s 68846 2128 68874 2184 4 bl_108
port 38 nsew
rlabel metal1 s 69310 2128 69338 2184 4 br_108
port 39 nsew
rlabel metal1 s 69906 2128 69934 2184 4 bl_109
port 40 nsew
rlabel metal1 s 69442 2128 69470 2184 4 br_109
port 41 nsew
rlabel metal1 s 70094 2128 70122 2184 4 bl_110
port 42 nsew
rlabel metal1 s 70558 2128 70586 2184 4 br_110
port 43 nsew
rlabel metal1 s 71154 2128 71182 2184 4 bl_111
port 44 nsew
rlabel metal1 s 70690 2128 70718 2184 4 br_111
port 45 nsew
rlabel metal1 s 71342 2128 71370 2184 4 bl_112
port 46 nsew
rlabel metal1 s 71806 2128 71834 2184 4 br_112
port 47 nsew
rlabel metal1 s 72402 2128 72430 2184 4 bl_113
port 48 nsew
rlabel metal1 s 71938 2128 71966 2184 4 br_113
port 49 nsew
rlabel metal1 s 72590 2128 72618 2184 4 bl_114
port 50 nsew
rlabel metal1 s 73054 2128 73082 2184 4 br_114
port 51 nsew
rlabel metal1 s 73650 2128 73678 2184 4 bl_115
port 52 nsew
rlabel metal1 s 73186 2128 73214 2184 4 br_115
port 53 nsew
rlabel metal1 s 73838 2128 73866 2184 4 bl_116
port 54 nsew
rlabel metal1 s 74302 2128 74330 2184 4 br_116
port 55 nsew
rlabel metal1 s 74898 2128 74926 2184 4 bl_117
port 56 nsew
rlabel metal1 s 74434 2128 74462 2184 4 br_117
port 57 nsew
rlabel metal1 s 75086 2128 75114 2184 4 bl_118
port 58 nsew
rlabel metal1 s 75550 2128 75578 2184 4 br_118
port 59 nsew
rlabel metal1 s 76146 2128 76174 2184 4 bl_119
port 60 nsew
rlabel metal1 s 75682 2128 75710 2184 4 br_119
port 61 nsew
rlabel metal1 s 76334 2128 76362 2184 4 bl_120
port 62 nsew
rlabel metal1 s 76798 2128 76826 2184 4 br_120
port 63 nsew
rlabel metal1 s 77394 2128 77422 2184 4 bl_121
port 64 nsew
rlabel metal1 s 76930 2128 76958 2184 4 br_121
port 65 nsew
rlabel metal1 s 77582 2128 77610 2184 4 bl_122
port 66 nsew
rlabel metal1 s 78046 2128 78074 2184 4 br_122
port 67 nsew
rlabel metal1 s 78642 2128 78670 2184 4 bl_123
port 68 nsew
rlabel metal1 s 78178 2128 78206 2184 4 br_123
port 69 nsew
rlabel metal1 s 78830 2128 78858 2184 4 bl_124
port 70 nsew
rlabel metal1 s 79294 2128 79322 2184 4 br_124
port 71 nsew
rlabel metal1 s 79890 2128 79918 2184 4 bl_125
port 72 nsew
rlabel metal1 s 79426 2128 79454 2184 4 br_125
port 73 nsew
rlabel metal1 s 80078 2128 80106 2184 4 bl_126
port 74 nsew
rlabel metal1 s 80542 2128 80570 2184 4 br_126
port 75 nsew
rlabel metal1 s 81138 2128 81166 2184 4 bl_127
port 76 nsew
rlabel metal1 s 80674 2128 80702 2184 4 br_127
port 77 nsew
rlabel metal1 s 58862 2128 58890 2184 4 bl_92
port 78 nsew
rlabel metal1 s 59326 2128 59354 2184 4 br_92
port 79 nsew
rlabel metal1 s 59922 2128 59950 2184 4 bl_93
port 80 nsew
rlabel metal1 s 59458 2128 59486 2184 4 br_93
port 81 nsew
rlabel metal1 s 60110 2128 60138 2184 4 bl_94
port 82 nsew
rlabel metal1 s 60574 2128 60602 2184 4 br_94
port 83 nsew
rlabel metal1 s 61170 2128 61198 2184 4 bl_95
port 84 nsew
rlabel metal1 s 60706 2128 60734 2184 4 br_95
port 85 nsew
rlabel metal1 s 41390 248 41418 868 4 bl_out_16
port 86 nsew
rlabel metal1 s 43886 248 43914 868 4 bl_out_17
port 87 nsew
rlabel metal1 s 46382 248 46410 868 4 bl_out_18
port 88 nsew
rlabel metal1 s 48878 248 48906 868 4 bl_out_19
port 89 nsew
rlabel metal1 s 51374 248 51402 868 4 bl_out_20
port 90 nsew
rlabel metal1 s 53870 248 53898 868 4 bl_out_21
port 91 nsew
rlabel metal1 s 56366 248 56394 868 4 bl_out_22
port 92 nsew
rlabel metal1 s 58862 248 58890 868 4 bl_out_23
port 93 nsew
rlabel metal1 s 41390 2128 41418 2184 4 bl_64
port 94 nsew
rlabel metal1 s 41854 2128 41882 2184 4 br_64
port 95 nsew
rlabel metal1 s 42450 2128 42478 2184 4 bl_65
port 96 nsew
rlabel metal1 s 41986 2128 42014 2184 4 br_65
port 97 nsew
rlabel metal1 s 42638 2128 42666 2184 4 bl_66
port 98 nsew
rlabel metal1 s 43102 2128 43130 2184 4 br_66
port 99 nsew
rlabel metal1 s 43698 2128 43726 2184 4 bl_67
port 100 nsew
rlabel metal1 s 43234 2128 43262 2184 4 br_67
port 101 nsew
rlabel metal1 s 43886 2128 43914 2184 4 bl_68
port 102 nsew
rlabel metal1 s 44350 2128 44378 2184 4 br_68
port 103 nsew
rlabel metal1 s 44946 2128 44974 2184 4 bl_69
port 104 nsew
rlabel metal1 s 44482 2128 44510 2184 4 br_69
port 105 nsew
rlabel metal1 s 45134 2128 45162 2184 4 bl_70
port 106 nsew
rlabel metal1 s 45598 2128 45626 2184 4 br_70
port 107 nsew
rlabel metal1 s 46194 2128 46222 2184 4 bl_71
port 108 nsew
rlabel metal1 s 45730 2128 45758 2184 4 br_71
port 109 nsew
rlabel metal1 s 46382 2128 46410 2184 4 bl_72
port 110 nsew
rlabel metal1 s 46846 2128 46874 2184 4 br_72
port 111 nsew
rlabel metal1 s 47442 2128 47470 2184 4 bl_73
port 112 nsew
rlabel metal1 s 46978 2128 47006 2184 4 br_73
port 113 nsew
rlabel metal1 s 47630 2128 47658 2184 4 bl_74
port 114 nsew
rlabel metal1 s 48094 2128 48122 2184 4 br_74
port 115 nsew
rlabel metal1 s 48690 2128 48718 2184 4 bl_75
port 116 nsew
rlabel metal1 s 48226 2128 48254 2184 4 br_75
port 117 nsew
rlabel metal1 s 48878 2128 48906 2184 4 bl_76
port 118 nsew
rlabel metal1 s 49342 2128 49370 2184 4 br_76
port 119 nsew
rlabel metal1 s 49938 2128 49966 2184 4 bl_77
port 120 nsew
rlabel metal1 s 49474 2128 49502 2184 4 br_77
port 121 nsew
rlabel metal1 s 50126 2128 50154 2184 4 bl_78
port 122 nsew
rlabel metal1 s 50590 2128 50618 2184 4 br_78
port 123 nsew
rlabel metal1 s 51186 2128 51214 2184 4 bl_79
port 124 nsew
rlabel metal1 s 50722 2128 50750 2184 4 br_79
port 125 nsew
rlabel metal1 s 51374 2128 51402 2184 4 bl_80
port 126 nsew
rlabel metal1 s 51838 2128 51866 2184 4 br_80
port 127 nsew
rlabel metal1 s 52434 2128 52462 2184 4 bl_81
port 128 nsew
rlabel metal1 s 51970 2128 51998 2184 4 br_81
port 129 nsew
rlabel metal1 s 52622 2128 52650 2184 4 bl_82
port 130 nsew
rlabel metal1 s 53086 2128 53114 2184 4 br_82
port 131 nsew
rlabel metal1 s 53682 2128 53710 2184 4 bl_83
port 132 nsew
rlabel metal1 s 53218 2128 53246 2184 4 br_83
port 133 nsew
rlabel metal1 s 53870 2128 53898 2184 4 bl_84
port 134 nsew
rlabel metal1 s 54334 2128 54362 2184 4 br_84
port 135 nsew
rlabel metal1 s 54930 2128 54958 2184 4 bl_85
port 136 nsew
rlabel metal1 s 54466 2128 54494 2184 4 br_85
port 137 nsew
rlabel metal1 s 55118 2128 55146 2184 4 bl_86
port 138 nsew
rlabel metal1 s 55582 2128 55610 2184 4 br_86
port 139 nsew
rlabel metal1 s 56178 2128 56206 2184 4 bl_87
port 140 nsew
rlabel metal1 s 55714 2128 55742 2184 4 br_87
port 141 nsew
rlabel metal1 s 56366 2128 56394 2184 4 bl_88
port 142 nsew
rlabel metal1 s 56830 2128 56858 2184 4 br_88
port 143 nsew
rlabel metal1 s 57426 2128 57454 2184 4 bl_89
port 144 nsew
rlabel metal1 s 56962 2128 56990 2184 4 br_89
port 145 nsew
rlabel metal1 s 57614 2128 57642 2184 4 bl_90
port 146 nsew
rlabel metal1 s 58078 2128 58106 2184 4 br_90
port 147 nsew
rlabel metal1 s 58674 2128 58702 2184 4 bl_91
port 148 nsew
rlabel metal1 s 58210 2128 58238 2184 4 br_91
port 149 nsew
rlabel metal1 s 36398 2128 36426 2184 4 bl_56
port 150 nsew
rlabel metal1 s 36862 2128 36890 2184 4 br_56
port 151 nsew
rlabel metal1 s 37458 2128 37486 2184 4 bl_57
port 152 nsew
rlabel metal1 s 36994 2128 37022 2184 4 br_57
port 153 nsew
rlabel metal1 s 37646 2128 37674 2184 4 bl_58
port 154 nsew
rlabel metal1 s 38110 2128 38138 2184 4 br_58
port 155 nsew
rlabel metal1 s 38706 2128 38734 2184 4 bl_59
port 156 nsew
rlabel metal1 s 38242 2128 38270 2184 4 br_59
port 157 nsew
rlabel metal1 s 38894 2128 38922 2184 4 bl_60
port 158 nsew
rlabel metal1 s 39358 2128 39386 2184 4 br_60
port 159 nsew
rlabel metal1 s 39954 2128 39982 2184 4 bl_61
port 160 nsew
rlabel metal1 s 39490 2128 39518 2184 4 br_61
port 161 nsew
rlabel metal1 s 40142 2128 40170 2184 4 bl_62
port 162 nsew
rlabel metal1 s 40606 2128 40634 2184 4 br_62
port 163 nsew
rlabel metal1 s 41202 2128 41230 2184 4 bl_63
port 164 nsew
rlabel metal1 s 40738 2128 40766 2184 4 br_63
port 165 nsew
rlabel metal1 s 21422 248 21450 868 4 bl_out_8
port 166 nsew
rlabel metal1 s 23918 248 23946 868 4 bl_out_9
port 167 nsew
rlabel metal1 s 26414 248 26442 868 4 bl_out_10
port 168 nsew
rlabel metal1 s 28910 248 28938 868 4 bl_out_11
port 169 nsew
rlabel metal1 s 31406 248 31434 868 4 bl_out_12
port 170 nsew
rlabel metal1 s 33902 248 33930 868 4 bl_out_13
port 171 nsew
rlabel metal1 s 36398 248 36426 868 4 bl_out_14
port 172 nsew
rlabel metal1 s 38894 248 38922 868 4 bl_out_15
port 173 nsew
rlabel metal1 s 21422 2128 21450 2184 4 bl_32
port 174 nsew
rlabel metal1 s 21886 2128 21914 2184 4 br_32
port 175 nsew
rlabel metal1 s 22482 2128 22510 2184 4 bl_33
port 176 nsew
rlabel metal1 s 22018 2128 22046 2184 4 br_33
port 177 nsew
rlabel metal1 s 22670 2128 22698 2184 4 bl_34
port 178 nsew
rlabel metal1 s 23134 2128 23162 2184 4 br_34
port 179 nsew
rlabel metal1 s 23730 2128 23758 2184 4 bl_35
port 180 nsew
rlabel metal1 s 23266 2128 23294 2184 4 br_35
port 181 nsew
rlabel metal1 s 23918 2128 23946 2184 4 bl_36
port 182 nsew
rlabel metal1 s 24382 2128 24410 2184 4 br_36
port 183 nsew
rlabel metal1 s 24978 2128 25006 2184 4 bl_37
port 184 nsew
rlabel metal1 s 24514 2128 24542 2184 4 br_37
port 185 nsew
rlabel metal1 s 25166 2128 25194 2184 4 bl_38
port 186 nsew
rlabel metal1 s 25630 2128 25658 2184 4 br_38
port 187 nsew
rlabel metal1 s 26226 2128 26254 2184 4 bl_39
port 188 nsew
rlabel metal1 s 25762 2128 25790 2184 4 br_39
port 189 nsew
rlabel metal1 s 26414 2128 26442 2184 4 bl_40
port 190 nsew
rlabel metal1 s 26878 2128 26906 2184 4 br_40
port 191 nsew
rlabel metal1 s 27474 2128 27502 2184 4 bl_41
port 192 nsew
rlabel metal1 s 27010 2128 27038 2184 4 br_41
port 193 nsew
rlabel metal1 s 27662 2128 27690 2184 4 bl_42
port 194 nsew
rlabel metal1 s 28126 2128 28154 2184 4 br_42
port 195 nsew
rlabel metal1 s 28722 2128 28750 2184 4 bl_43
port 196 nsew
rlabel metal1 s 28258 2128 28286 2184 4 br_43
port 197 nsew
rlabel metal1 s 28910 2128 28938 2184 4 bl_44
port 198 nsew
rlabel metal1 s 29374 2128 29402 2184 4 br_44
port 199 nsew
rlabel metal1 s 29970 2128 29998 2184 4 bl_45
port 200 nsew
rlabel metal1 s 29506 2128 29534 2184 4 br_45
port 201 nsew
rlabel metal1 s 30158 2128 30186 2184 4 bl_46
port 202 nsew
rlabel metal1 s 30622 2128 30650 2184 4 br_46
port 203 nsew
rlabel metal1 s 31218 2128 31246 2184 4 bl_47
port 204 nsew
rlabel metal1 s 30754 2128 30782 2184 4 br_47
port 205 nsew
rlabel metal1 s 31406 2128 31434 2184 4 bl_48
port 206 nsew
rlabel metal1 s 31870 2128 31898 2184 4 br_48
port 207 nsew
rlabel metal1 s 32466 2128 32494 2184 4 bl_49
port 208 nsew
rlabel metal1 s 32002 2128 32030 2184 4 br_49
port 209 nsew
rlabel metal1 s 32654 2128 32682 2184 4 bl_50
port 210 nsew
rlabel metal1 s 33118 2128 33146 2184 4 br_50
port 211 nsew
rlabel metal1 s 33714 2128 33742 2184 4 bl_51
port 212 nsew
rlabel metal1 s 33250 2128 33278 2184 4 br_51
port 213 nsew
rlabel metal1 s 33902 2128 33930 2184 4 bl_52
port 214 nsew
rlabel metal1 s 34366 2128 34394 2184 4 br_52
port 215 nsew
rlabel metal1 s 34962 2128 34990 2184 4 bl_53
port 216 nsew
rlabel metal1 s 34498 2128 34526 2184 4 br_53
port 217 nsew
rlabel metal1 s 35150 2128 35178 2184 4 bl_54
port 218 nsew
rlabel metal1 s 35614 2128 35642 2184 4 br_54
port 219 nsew
rlabel metal1 s 36210 2128 36238 2184 4 bl_55
port 220 nsew
rlabel metal1 s 35746 2128 35774 2184 4 br_55
port 221 nsew
rlabel metal1 s 13934 2128 13962 2184 4 bl_20
port 222 nsew
rlabel metal1 s 14398 2128 14426 2184 4 br_20
port 223 nsew
rlabel metal1 s 14994 2128 15022 2184 4 bl_21
port 224 nsew
rlabel metal1 s 14530 2128 14558 2184 4 br_21
port 225 nsew
rlabel metal1 s 15182 2128 15210 2184 4 bl_22
port 226 nsew
rlabel metal1 s 15646 2128 15674 2184 4 br_22
port 227 nsew
rlabel metal1 s 16242 2128 16270 2184 4 bl_23
port 228 nsew
rlabel metal1 s 15778 2128 15806 2184 4 br_23
port 229 nsew
rlabel metal1 s 16430 2128 16458 2184 4 bl_24
port 230 nsew
rlabel metal1 s 16894 2128 16922 2184 4 br_24
port 231 nsew
rlabel metal1 s 17490 2128 17518 2184 4 bl_25
port 232 nsew
rlabel metal1 s 17026 2128 17054 2184 4 br_25
port 233 nsew
rlabel metal1 s 17678 2128 17706 2184 4 bl_26
port 234 nsew
rlabel metal1 s 18142 2128 18170 2184 4 br_26
port 235 nsew
rlabel metal1 s 18738 2128 18766 2184 4 bl_27
port 236 nsew
rlabel metal1 s 18274 2128 18302 2184 4 br_27
port 237 nsew
rlabel metal1 s 18926 2128 18954 2184 4 bl_28
port 238 nsew
rlabel metal1 s 19390 2128 19418 2184 4 br_28
port 239 nsew
rlabel metal1 s 19986 2128 20014 2184 4 bl_29
port 240 nsew
rlabel metal1 s 19522 2128 19550 2184 4 br_29
port 241 nsew
rlabel metal1 s 20174 2128 20202 2184 4 bl_30
port 242 nsew
rlabel metal1 s 20638 2128 20666 2184 4 br_30
port 243 nsew
rlabel metal1 s 21234 2128 21262 2184 4 bl_31
port 244 nsew
rlabel metal1 s 20770 2128 20798 2184 4 br_31
port 245 nsew
rlabel metal1 s 1454 248 1482 868 4 bl_out_0
port 246 nsew
rlabel metal1 s 3950 248 3978 868 4 bl_out_1
port 247 nsew
rlabel metal1 s 6446 248 6474 868 4 bl_out_2
port 248 nsew
rlabel metal1 s 8942 248 8970 868 4 bl_out_3
port 249 nsew
rlabel metal1 s 11438 248 11466 868 4 bl_out_4
port 250 nsew
rlabel metal1 s 13934 248 13962 868 4 bl_out_5
port 251 nsew
rlabel metal1 s 16430 248 16458 868 4 bl_out_6
port 252 nsew
rlabel metal1 s 18926 248 18954 868 4 bl_out_7
port 253 nsew
rlabel metal1 s 1454 2128 1482 2184 4 bl_0
port 254 nsew
rlabel metal1 s 1918 2128 1946 2184 4 br_0
port 255 nsew
rlabel metal1 s 2514 2128 2542 2184 4 bl_1
port 256 nsew
rlabel metal1 s 2050 2128 2078 2184 4 br_1
port 257 nsew
rlabel metal1 s 2702 2128 2730 2184 4 bl_2
port 258 nsew
rlabel metal1 s 3166 2128 3194 2184 4 br_2
port 259 nsew
rlabel metal1 s 3762 2128 3790 2184 4 bl_3
port 260 nsew
rlabel metal1 s 3298 2128 3326 2184 4 br_3
port 261 nsew
rlabel metal1 s 3950 2128 3978 2184 4 bl_4
port 262 nsew
rlabel metal1 s 4414 2128 4442 2184 4 br_4
port 263 nsew
rlabel metal1 s 5010 2128 5038 2184 4 bl_5
port 264 nsew
rlabel metal1 s 4546 2128 4574 2184 4 br_5
port 265 nsew
rlabel metal1 s 5198 2128 5226 2184 4 bl_6
port 266 nsew
rlabel metal1 s 5662 2128 5690 2184 4 br_6
port 267 nsew
rlabel metal1 s 6258 2128 6286 2184 4 bl_7
port 268 nsew
rlabel metal1 s 5794 2128 5822 2184 4 br_7
port 269 nsew
rlabel metal1 s 6446 2128 6474 2184 4 bl_8
port 270 nsew
rlabel metal1 s 6910 2128 6938 2184 4 br_8
port 271 nsew
rlabel metal1 s 7506 2128 7534 2184 4 bl_9
port 272 nsew
rlabel metal1 s 7042 2128 7070 2184 4 br_9
port 273 nsew
rlabel metal1 s 7694 2128 7722 2184 4 bl_10
port 274 nsew
rlabel metal1 s 8158 2128 8186 2184 4 br_10
port 275 nsew
rlabel metal1 s 8754 2128 8782 2184 4 bl_11
port 276 nsew
rlabel metal1 s 8290 2128 8318 2184 4 br_11
port 277 nsew
rlabel metal1 s 8942 2128 8970 2184 4 bl_12
port 278 nsew
rlabel metal1 s 9406 2128 9434 2184 4 br_12
port 279 nsew
rlabel metal1 s 10002 2128 10030 2184 4 bl_13
port 280 nsew
rlabel metal1 s 9538 2128 9566 2184 4 br_13
port 281 nsew
rlabel metal1 s 10190 2128 10218 2184 4 bl_14
port 282 nsew
rlabel metal1 s 10654 2128 10682 2184 4 br_14
port 283 nsew
rlabel metal1 s 11250 2128 11278 2184 4 bl_15
port 284 nsew
rlabel metal1 s 10786 2128 10814 2184 4 br_15
port 285 nsew
rlabel metal1 s 11438 2128 11466 2184 4 bl_16
port 286 nsew
rlabel metal1 s 11902 2128 11930 2184 4 br_16
port 287 nsew
rlabel metal1 s 12498 2128 12526 2184 4 bl_17
port 288 nsew
rlabel metal1 s 12034 2128 12062 2184 4 br_17
port 289 nsew
rlabel metal1 s 12686 2128 12714 2184 4 bl_18
port 290 nsew
rlabel metal1 s 13150 2128 13178 2184 4 br_18
port 291 nsew
rlabel metal1 s 13746 2128 13774 2184 4 bl_19
port 292 nsew
rlabel metal1 s 13282 2128 13310 2184 4 br_19
port 293 nsew
rlabel metal1 s 1918 124 1946 868 4 br_out_0
port 294 nsew
rlabel metal1 s 21886 124 21914 868 4 br_out_8
port 295 nsew
rlabel metal1 s 11902 124 11930 868 4 br_out_4
port 296 nsew
rlabel metal1 s 24382 124 24410 868 4 br_out_9
port 297 nsew
rlabel metal1 s 6910 124 6938 868 4 br_out_2
port 298 nsew
rlabel metal1 s 26878 124 26906 868 4 br_out_10
port 299 nsew
rlabel metal1 s 14398 124 14426 868 4 br_out_5
port 300 nsew
rlabel metal1 s 29374 124 29402 868 4 br_out_11
port 301 nsew
rlabel metal1 s 4414 124 4442 868 4 br_out_1
port 302 nsew
rlabel metal1 s 31870 124 31898 868 4 br_out_12
port 303 nsew
rlabel metal1 s 16894 124 16922 868 4 br_out_6
port 304 nsew
rlabel metal1 s 34366 124 34394 868 4 br_out_13
port 305 nsew
rlabel metal1 s 9406 124 9434 868 4 br_out_3
port 306 nsew
rlabel metal1 s 36862 124 36890 868 4 br_out_14
port 307 nsew
rlabel metal1 s 19390 124 19418 868 4 br_out_7
port 308 nsew
rlabel metal1 s 39358 124 39386 868 4 br_out_15
port 309 nsew
rlabel metal1 s 41854 124 41882 868 4 br_out_16
port 310 nsew
rlabel metal1 s 61822 124 61850 868 4 br_out_24
port 311 nsew
rlabel metal1 s 51838 124 51866 868 4 br_out_20
port 312 nsew
rlabel metal1 s 64318 124 64346 868 4 br_out_25
port 313 nsew
rlabel metal1 s 46846 124 46874 868 4 br_out_18
port 314 nsew
rlabel metal1 s 66814 124 66842 868 4 br_out_26
port 315 nsew
rlabel metal1 s 54334 124 54362 868 4 br_out_21
port 316 nsew
rlabel metal1 s 69310 124 69338 868 4 br_out_27
port 317 nsew
rlabel metal1 s 44350 124 44378 868 4 br_out_17
port 318 nsew
rlabel metal1 s 71806 124 71834 868 4 br_out_28
port 319 nsew
rlabel metal1 s 56830 124 56858 868 4 br_out_22
port 320 nsew
rlabel metal1 s 74302 124 74330 868 4 br_out_29
port 321 nsew
rlabel metal1 s 49342 124 49370 868 4 br_out_19
port 322 nsew
rlabel metal1 s 76798 124 76826 868 4 br_out_30
port 323 nsew
rlabel metal1 s 59326 124 59354 868 4 br_out_23
port 324 nsew
rlabel metal1 s 79294 124 79322 868 4 br_out_31
port 325 nsew
<< properties >>
string FIXED_BBOX 80655 87 80721 161
string GDS_END 1357146
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 1142012
<< end >>
