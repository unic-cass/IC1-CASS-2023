magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 1011 203
rect 30 -17 64 21
<< locali >>
rect 543 451 995 485
rect 950 357 995 451
rect 86 199 156 265
rect 494 215 712 255
rect 862 199 927 323
rect 116 145 156 199
rect 961 93 995 357
rect 543 59 995 93
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 427 69 493
rect 103 451 169 527
rect 271 451 337 527
rect 371 427 416 493
rect 455 435 505 527
rect 17 333 52 427
rect 382 401 416 427
rect 543 401 870 417
rect 187 367 347 401
rect 382 383 870 401
rect 382 367 577 383
rect 313 333 347 367
rect 627 333 693 343
rect 17 299 279 333
rect 313 299 693 333
rect 17 135 52 299
rect 245 265 279 299
rect 245 231 397 265
rect 331 215 397 231
rect 17 69 69 135
rect 203 115 251 187
rect 103 17 167 109
rect 287 17 337 177
rect 371 147 693 181
rect 371 59 405 147
rect 627 131 693 147
rect 770 165 821 187
rect 770 131 869 165
rect 455 17 489 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< obsm1 >>
rect 202 184 260 193
rect 758 184 816 193
rect 202 156 816 184
rect 202 147 260 156
rect 758 147 816 156
<< labels >>
rlabel locali s 494 215 712 255 6 A0
port 1 nsew signal input
rlabel locali s 862 199 927 323 6 A1
port 2 nsew signal input
rlabel locali s 116 145 156 199 6 S
port 3 nsew signal input
rlabel locali s 86 199 156 265 6 S
port 3 nsew signal input
rlabel metal1 s 0 -48 1012 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1011 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 543 59 995 93 6 Y
port 8 nsew signal output
rlabel locali s 961 93 995 357 6 Y
port 8 nsew signal output
rlabel locali s 950 357 995 451 6 Y
port 8 nsew signal output
rlabel locali s 543 451 995 485 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1705622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1697608
<< end >>
