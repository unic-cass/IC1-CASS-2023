magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 10 43 764 289
rect -26 -43 794 43
<< mvnmos >>
rect 93 113 193 263
rect 249 113 349 263
rect 405 113 505 263
rect 581 113 681 263
<< mvpmos >>
rect 107 443 207 743
rect 249 443 349 743
rect 420 443 520 743
rect 562 443 662 743
<< mvndiff >>
rect 36 255 93 263
rect 36 221 48 255
rect 82 221 93 255
rect 36 155 93 221
rect 36 121 48 155
rect 82 121 93 155
rect 36 113 93 121
rect 193 255 249 263
rect 193 221 204 255
rect 238 221 249 255
rect 193 157 249 221
rect 193 123 204 157
rect 238 123 249 157
rect 193 113 249 123
rect 349 255 405 263
rect 349 221 360 255
rect 394 221 405 255
rect 349 155 405 221
rect 349 121 360 155
rect 394 121 405 155
rect 349 113 405 121
rect 505 255 581 263
rect 505 221 516 255
rect 550 221 581 255
rect 505 155 581 221
rect 505 121 516 155
rect 550 121 581 155
rect 505 113 581 121
rect 681 255 738 263
rect 681 221 692 255
rect 726 221 738 255
rect 681 155 738 221
rect 681 121 692 155
rect 726 121 738 155
rect 681 113 738 121
<< mvpdiff >>
rect 50 735 107 743
rect 50 701 62 735
rect 96 701 107 735
rect 50 654 107 701
rect 50 620 62 654
rect 96 620 107 654
rect 50 571 107 620
rect 50 537 62 571
rect 96 537 107 571
rect 50 490 107 537
rect 50 456 62 490
rect 96 456 107 490
rect 50 443 107 456
rect 207 443 249 743
rect 349 735 420 743
rect 349 701 375 735
rect 409 701 420 735
rect 349 652 420 701
rect 349 618 375 652
rect 409 618 420 652
rect 349 568 420 618
rect 349 534 375 568
rect 409 534 420 568
rect 349 485 420 534
rect 349 451 375 485
rect 409 451 420 485
rect 349 443 420 451
rect 520 443 562 743
rect 662 735 719 743
rect 662 701 673 735
rect 707 701 719 735
rect 662 655 719 701
rect 662 621 673 655
rect 707 621 719 655
rect 662 574 719 621
rect 662 540 673 574
rect 707 540 719 574
rect 662 494 719 540
rect 662 460 673 494
rect 707 460 719 494
rect 662 443 719 460
<< mvndiffc >>
rect 48 221 82 255
rect 48 121 82 155
rect 204 221 238 255
rect 204 123 238 157
rect 360 221 394 255
rect 360 121 394 155
rect 516 221 550 255
rect 516 121 550 155
rect 692 221 726 255
rect 692 121 726 155
<< mvpdiffc >>
rect 62 701 96 735
rect 62 620 96 654
rect 62 537 96 571
rect 62 456 96 490
rect 375 701 409 735
rect 375 618 409 652
rect 375 534 409 568
rect 375 451 409 485
rect 673 701 707 735
rect 673 621 707 655
rect 673 540 707 574
rect 673 460 707 494
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
<< poly >>
rect 107 743 207 769
rect 249 743 349 769
rect 420 743 520 769
rect 562 743 662 769
rect 107 385 207 443
rect 40 357 207 385
rect 40 323 60 357
rect 94 323 207 357
rect 40 285 207 323
rect 249 346 349 443
rect 420 421 520 443
rect 249 312 269 346
rect 303 312 349 346
rect 93 263 193 285
rect 249 263 349 312
rect 405 395 520 421
rect 405 361 466 395
rect 500 361 520 395
rect 405 321 520 361
rect 562 417 662 443
rect 562 395 681 417
rect 562 361 625 395
rect 659 361 681 395
rect 405 263 505 321
rect 562 289 681 361
rect 581 263 681 289
rect 93 87 193 113
rect 249 87 349 113
rect 405 87 505 113
rect 581 87 681 113
<< polycont >>
rect 60 323 94 357
rect 269 312 303 346
rect 466 361 500 395
rect 625 361 659 395
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 18 735 269 751
rect 18 701 19 735
rect 53 701 62 735
rect 125 701 163 735
rect 197 701 235 735
rect 18 654 269 701
rect 18 620 62 654
rect 96 620 269 654
rect 375 735 409 751
rect 375 652 409 701
rect 18 571 269 620
rect 18 537 62 571
rect 96 537 269 571
rect 18 490 269 537
rect 18 456 62 490
rect 96 456 269 490
rect 305 618 375 652
rect 305 568 409 618
rect 305 534 375 568
rect 305 485 409 534
rect 305 451 375 485
rect 461 735 723 751
rect 461 701 467 735
rect 501 701 539 735
rect 573 701 611 735
rect 645 701 673 735
rect 717 701 723 735
rect 461 655 723 701
rect 461 621 673 655
rect 707 621 723 655
rect 461 574 723 621
rect 461 540 673 574
rect 707 540 723 574
rect 461 494 723 540
rect 461 460 673 494
rect 707 460 723 494
rect 305 435 409 451
rect 305 420 359 435
rect 147 386 359 420
rect 450 395 551 424
rect 25 357 110 373
rect 25 323 60 357
rect 94 323 110 357
rect 25 307 110 323
rect 147 271 181 386
rect 450 361 466 395
rect 500 361 551 395
rect 601 395 743 424
rect 601 361 625 395
rect 659 361 743 395
rect 217 346 319 350
rect 217 312 269 346
rect 303 312 319 346
rect 217 307 319 312
rect 360 291 734 325
rect 32 255 98 271
rect 32 221 48 255
rect 82 221 98 255
rect 32 155 98 221
rect 32 121 48 155
rect 82 121 98 155
rect 147 255 254 271
rect 147 221 204 255
rect 238 221 254 255
rect 147 157 254 221
rect 147 123 204 157
rect 238 123 254 157
rect 360 255 394 291
rect 684 255 734 291
rect 360 155 394 221
rect 32 87 98 121
rect 360 87 394 121
rect 32 53 394 87
rect 430 221 516 255
rect 550 221 650 255
rect 430 155 650 221
rect 430 121 516 155
rect 550 121 650 155
rect 430 113 650 121
rect 430 79 440 113
rect 474 79 512 113
rect 546 79 584 113
rect 618 79 650 113
rect 684 221 692 255
rect 726 221 734 255
rect 684 155 734 221
rect 684 121 692 155
rect 726 121 734 155
rect 684 105 734 121
rect 430 73 650 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 19 701 53 735
rect 91 701 96 735
rect 96 701 125 735
rect 163 701 197 735
rect 235 701 269 735
rect 467 701 501 735
rect 539 701 573 735
rect 611 701 645 735
rect 683 701 707 735
rect 707 701 717 735
rect 440 79 474 113
rect 512 79 546 113
rect 584 79 618 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 19 735
rect 53 701 91 735
rect 125 701 163 735
rect 197 701 235 735
rect 269 701 467 735
rect 501 701 539 735
rect 573 701 611 735
rect 645 701 683 735
rect 717 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 440 113
rect 474 79 512 113
rect 546 79 584 113
rect 618 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o22ai_1
flabel metal1 s 0 51 768 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 768 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 768 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 768 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 612 353 646 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 768 814
string GDS_END 386136
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 376348
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
