magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 5 21 735 203
rect 29 -17 63 21
rect 395 -13 429 21
<< locali >>
rect 29 176 106 492
rect 157 210 247 491
rect 287 210 354 491
rect 388 280 443 491
rect 388 210 454 280
rect 488 199 545 280
rect 581 204 708 258
rect 29 163 460 176
rect 29 141 484 163
rect 29 140 275 141
rect 209 52 275 140
rect 418 61 484 141
rect 581 70 618 204
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 479 350 525 492
rect 560 384 626 527
rect 662 350 701 492
rect 479 316 701 350
rect 63 17 126 105
rect 310 17 376 107
rect 654 17 702 152
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 488 199 545 280 6 A1
port 1 nsew signal input
rlabel locali s 581 70 618 204 6 A2
port 2 nsew signal input
rlabel locali s 581 204 708 258 6 A2
port 2 nsew signal input
rlabel locali s 388 210 454 280 6 B1
port 3 nsew signal input
rlabel locali s 388 280 443 491 6 B1
port 3 nsew signal input
rlabel locali s 287 210 354 491 6 C1
port 4 nsew signal input
rlabel locali s 157 210 247 491 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 395 -13 429 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 5 21 735 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 418 61 484 141 6 Y
port 10 nsew signal output
rlabel locali s 209 52 275 140 6 Y
port 10 nsew signal output
rlabel locali s 29 140 275 141 6 Y
port 10 nsew signal output
rlabel locali s 29 141 484 163 6 Y
port 10 nsew signal output
rlabel locali s 29 163 460 176 6 Y
port 10 nsew signal output
rlabel locali s 29 176 106 492 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3798426
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3790644
<< end >>
