magic
tech sky130B
timestamp 1676037725
<< obsli1 >>
rect 0 693 27 738
rect 831 728 858 752
rect 44 711 858 728
rect 0 676 814 693
rect 0 623 27 676
rect 831 658 858 711
rect 44 641 858 658
rect 0 606 814 623
rect 0 553 27 606
rect 831 588 858 641
rect 44 571 858 588
rect 0 536 814 553
rect 0 483 27 536
rect 831 518 858 571
rect 44 501 858 518
rect 0 466 814 483
rect 0 413 27 466
rect 831 448 858 501
rect 44 431 858 448
rect 0 396 814 413
rect 0 343 27 396
rect 831 378 858 431
rect 44 361 858 378
rect 0 326 814 343
rect 0 273 27 326
rect 831 308 858 361
rect 44 291 858 308
rect 0 256 814 273
rect 0 203 27 256
rect 831 238 858 291
rect 44 221 858 238
rect 0 186 814 203
rect 0 133 27 186
rect 831 168 858 221
rect 44 151 858 168
rect 0 116 814 133
rect 0 63 27 116
rect 831 98 858 151
rect 44 81 858 98
rect 0 46 814 63
rect 831 46 858 81
rect 0 32 27 46
<< obsm1 >>
rect 0 752 858 784
rect 0 32 27 738
rect 44 32 58 738
rect 72 46 86 752
rect 100 32 114 738
rect 128 46 142 752
rect 156 32 170 738
rect 184 46 198 752
rect 212 32 226 738
rect 240 46 254 752
rect 268 32 282 738
rect 296 46 310 752
rect 324 32 338 738
rect 352 46 366 752
rect 380 32 394 738
rect 408 46 422 752
rect 436 32 450 738
rect 464 46 478 752
rect 492 32 506 738
rect 520 46 534 752
rect 548 32 562 738
rect 576 46 590 752
rect 604 32 618 738
rect 632 46 646 752
rect 660 32 674 738
rect 688 46 702 752
rect 716 32 730 738
rect 744 46 758 752
rect 772 32 786 738
rect 800 46 814 752
rect 831 46 858 752
rect 0 0 858 32
<< obsm2 >>
rect 0 752 858 784
rect 0 32 27 738
rect 44 46 58 752
rect 72 32 86 738
rect 100 46 114 752
rect 128 32 142 738
rect 156 46 170 752
rect 184 32 198 738
rect 212 46 226 752
rect 240 32 254 738
rect 268 46 282 752
rect 296 32 310 738
rect 324 46 338 752
rect 352 32 366 738
rect 380 46 394 752
rect 408 32 422 738
rect 436 46 450 752
rect 464 32 478 738
rect 492 46 506 752
rect 520 32 534 738
rect 548 46 562 752
rect 576 32 590 738
rect 604 46 618 752
rect 632 32 646 738
rect 660 46 674 752
rect 688 32 702 738
rect 716 46 730 752
rect 744 32 758 738
rect 772 46 786 752
rect 800 32 814 738
rect 831 46 858 752
rect 0 0 858 32
<< properties >>
string FIXED_BBOX 0 0 858 784
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 256840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 241220
<< end >>
