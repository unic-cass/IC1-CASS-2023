magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 15 67 627 203
rect 29 21 627 67
rect 29 -17 63 21
<< scnmos >>
rect 94 93 124 177
rect 202 47 232 177
rect 286 47 316 177
rect 393 47 423 177
rect 501 47 531 177
<< scpmoshvt >>
rect 105 297 135 381
rect 202 297 232 497
rect 286 297 316 497
rect 393 297 423 497
rect 501 297 531 497
<< ndiff >>
rect 41 139 94 177
rect 41 105 49 139
rect 83 105 94 139
rect 41 93 94 105
rect 124 93 202 177
rect 139 59 147 93
rect 181 59 202 93
rect 139 47 202 59
rect 232 47 286 177
rect 316 47 393 177
rect 423 47 501 177
rect 531 161 601 177
rect 531 127 555 161
rect 589 127 601 161
rect 531 93 601 127
rect 531 59 555 93
rect 589 59 601 93
rect 531 47 601 59
<< pdiff >>
rect 150 485 202 497
rect 150 451 158 485
rect 192 451 202 485
rect 150 417 202 451
rect 150 383 158 417
rect 192 383 202 417
rect 150 381 202 383
rect 53 369 105 381
rect 53 335 61 369
rect 95 335 105 369
rect 53 297 105 335
rect 135 349 202 381
rect 135 315 158 349
rect 192 315 202 349
rect 135 297 202 315
rect 232 485 286 497
rect 232 451 242 485
rect 276 451 286 485
rect 232 417 286 451
rect 232 383 242 417
rect 276 383 286 417
rect 232 349 286 383
rect 232 315 242 349
rect 276 315 286 349
rect 232 297 286 315
rect 316 485 393 497
rect 316 451 338 485
rect 372 451 393 485
rect 316 417 393 451
rect 316 383 338 417
rect 372 383 393 417
rect 316 297 393 383
rect 423 484 501 497
rect 423 450 433 484
rect 467 450 501 484
rect 423 416 501 450
rect 423 382 433 416
rect 467 382 501 416
rect 423 348 501 382
rect 423 314 433 348
rect 467 314 501 348
rect 423 297 501 314
rect 531 485 587 497
rect 531 451 541 485
rect 575 451 587 485
rect 531 417 587 451
rect 531 383 541 417
rect 575 383 587 417
rect 531 297 587 383
<< ndiffc >>
rect 49 105 83 139
rect 147 59 181 93
rect 555 127 589 161
rect 555 59 589 93
<< pdiffc >>
rect 158 451 192 485
rect 158 383 192 417
rect 61 335 95 369
rect 158 315 192 349
rect 242 451 276 485
rect 242 383 276 417
rect 242 315 276 349
rect 338 451 372 485
rect 338 383 372 417
rect 433 450 467 484
rect 433 382 467 416
rect 433 314 467 348
rect 541 451 575 485
rect 541 383 575 417
<< poly >>
rect 202 497 232 523
rect 286 497 316 523
rect 393 497 423 523
rect 501 497 531 523
rect 105 381 135 407
rect 105 265 135 297
rect 202 265 232 297
rect 286 265 316 297
rect 393 265 423 297
rect 501 265 531 297
rect 69 249 135 265
rect 69 215 85 249
rect 119 215 135 249
rect 69 199 135 215
rect 177 249 243 265
rect 177 215 193 249
rect 227 215 243 249
rect 177 199 243 215
rect 285 249 351 265
rect 285 215 301 249
rect 335 215 351 249
rect 285 199 351 215
rect 393 249 447 265
rect 393 215 403 249
rect 437 215 447 249
rect 393 199 447 215
rect 501 249 567 265
rect 501 215 517 249
rect 551 215 567 249
rect 501 199 567 215
rect 94 177 124 199
rect 202 177 232 199
rect 286 177 316 199
rect 393 177 423 199
rect 501 177 531 199
rect 94 67 124 93
rect 202 21 232 47
rect 286 21 316 47
rect 393 21 423 47
rect 501 21 531 47
<< polycont >>
rect 85 215 119 249
rect 193 215 227 249
rect 301 215 335 249
rect 403 215 437 249
rect 517 215 551 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 142 485 192 527
rect 142 451 158 485
rect 142 417 192 451
rect 17 369 102 385
rect 17 335 61 369
rect 95 335 102 369
rect 17 319 102 335
rect 142 383 158 417
rect 142 349 192 383
rect 17 165 51 319
rect 142 315 158 349
rect 142 299 192 315
rect 226 485 292 493
rect 226 451 242 485
rect 276 451 292 485
rect 226 417 292 451
rect 226 383 242 417
rect 276 383 292 417
rect 226 349 292 383
rect 326 485 383 527
rect 326 451 338 485
rect 372 451 383 485
rect 326 417 383 451
rect 326 383 338 417
rect 372 383 383 417
rect 326 367 383 383
rect 417 484 483 493
rect 417 450 433 484
rect 467 450 483 484
rect 417 416 483 450
rect 417 382 433 416
rect 467 382 483 416
rect 226 315 242 349
rect 276 333 292 349
rect 417 348 483 382
rect 541 485 584 527
rect 575 451 584 485
rect 541 417 584 451
rect 575 383 584 417
rect 541 367 584 383
rect 417 333 433 348
rect 276 315 433 333
rect 226 314 433 315
rect 467 333 483 348
rect 467 314 627 333
rect 226 299 627 314
rect 85 249 155 265
rect 119 215 155 249
rect 85 199 155 215
rect 193 249 247 265
rect 227 215 247 249
rect 193 199 247 215
rect 301 249 351 265
rect 335 215 351 249
rect 17 139 267 165
rect 301 153 351 215
rect 385 249 437 265
rect 385 215 403 249
rect 385 153 437 215
rect 471 249 551 265
rect 471 215 517 249
rect 471 199 551 215
rect 17 105 49 139
rect 83 131 267 139
rect 83 105 95 131
rect 17 89 95 105
rect 231 119 267 131
rect 471 119 505 199
rect 585 165 627 299
rect 131 93 197 97
rect 131 59 147 93
rect 181 59 197 93
rect 231 85 505 119
rect 539 161 627 165
rect 539 127 555 161
rect 589 127 627 161
rect 539 93 627 127
rect 131 17 197 59
rect 539 59 555 93
rect 589 59 627 93
rect 539 51 627 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 581 85 615 119 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 305 221 339 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand4b_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1900974
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1895160
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
