magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 26 3332 8008 3632
rect 26 3296 520 3332
tri 204 3280 220 3296 ne
rect 220 3160 520 3296
tri 520 3190 662 3332 nw
tri 902 3190 1044 3332 ne
rect 1044 3160 1344 3332
tri 1344 3190 1486 3332 nw
tri 1726 3190 1868 3332 ne
rect 1868 3160 2168 3332
tri 2168 3190 2310 3332 nw
tri 2550 3190 2692 3332 ne
rect 2692 3160 2992 3332
tri 2992 3190 3134 3332 nw
tri 3374 3190 3516 3332 ne
rect 3516 3160 3816 3332
tri 3816 3190 3958 3332 nw
tri 4488 3190 4630 3332 ne
rect 4630 3160 4930 3332
tri 4930 3190 5072 3332 nw
tri 5312 3190 5454 3332 ne
rect 5454 3160 5754 3332
tri 5754 3190 5896 3332 nw
tri 6136 3190 6278 3332 ne
rect 6278 3160 6578 3332
tri 6578 3190 6720 3332 nw
tri 6960 3190 7102 3332 ne
rect 7102 3160 7402 3332
tri 7402 3190 7544 3332 nw
tri 7784 3190 7926 3332 ne
rect 7926 3190 8008 3332
use sky130_fd_io__gnd2gnd_sub_dnwl  sky130_fd_io__gnd2gnd_sub_dnwl_0
timestamp 1676037725
transform 1 0 0 0 1 0
box 26 26 3956 3333
use sky130_fd_io__gnd2gnd_sub_dnwl  sky130_fd_io__gnd2gnd_sub_dnwl_1
timestamp 1676037725
transform -1 0 8034 0 1 0
box 26 26 3956 3333
<< properties >>
string GDS_END 8056168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8053780
<< end >>
