magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -54 284 4632 454
rect -59 116 4637 284
rect -54 -54 4632 116
<< scpmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
rect 384 0 414 400
rect 492 0 522 400
rect 600 0 630 400
rect 708 0 738 400
rect 816 0 846 400
rect 924 0 954 400
rect 1032 0 1062 400
rect 1140 0 1170 400
rect 1248 0 1278 400
rect 1356 0 1386 400
rect 1464 0 1494 400
rect 1572 0 1602 400
rect 1680 0 1710 400
rect 1788 0 1818 400
rect 1896 0 1926 400
rect 2004 0 2034 400
rect 2112 0 2142 400
rect 2220 0 2250 400
rect 2328 0 2358 400
rect 2436 0 2466 400
rect 2544 0 2574 400
rect 2652 0 2682 400
rect 2760 0 2790 400
rect 2868 0 2898 400
rect 2976 0 3006 400
rect 3084 0 3114 400
rect 3192 0 3222 400
rect 3300 0 3330 400
rect 3408 0 3438 400
rect 3516 0 3546 400
rect 3624 0 3654 400
rect 3732 0 3762 400
rect 3840 0 3870 400
rect 3948 0 3978 400
rect 4056 0 4086 400
rect 4164 0 4194 400
rect 4272 0 4302 400
rect 4380 0 4410 400
rect 4488 0 4518 400
<< pdiff >>
rect 0 217 60 400
rect 0 183 8 217
rect 42 183 60 217
rect 0 0 60 183
rect 90 217 168 400
rect 90 183 112 217
rect 146 183 168 217
rect 90 0 168 183
rect 198 217 276 400
rect 198 183 220 217
rect 254 183 276 217
rect 198 0 276 183
rect 306 217 384 400
rect 306 183 328 217
rect 362 183 384 217
rect 306 0 384 183
rect 414 217 492 400
rect 414 183 436 217
rect 470 183 492 217
rect 414 0 492 183
rect 522 217 600 400
rect 522 183 544 217
rect 578 183 600 217
rect 522 0 600 183
rect 630 217 708 400
rect 630 183 652 217
rect 686 183 708 217
rect 630 0 708 183
rect 738 217 816 400
rect 738 183 760 217
rect 794 183 816 217
rect 738 0 816 183
rect 846 217 924 400
rect 846 183 868 217
rect 902 183 924 217
rect 846 0 924 183
rect 954 217 1032 400
rect 954 183 976 217
rect 1010 183 1032 217
rect 954 0 1032 183
rect 1062 217 1140 400
rect 1062 183 1084 217
rect 1118 183 1140 217
rect 1062 0 1140 183
rect 1170 217 1248 400
rect 1170 183 1192 217
rect 1226 183 1248 217
rect 1170 0 1248 183
rect 1278 217 1356 400
rect 1278 183 1300 217
rect 1334 183 1356 217
rect 1278 0 1356 183
rect 1386 217 1464 400
rect 1386 183 1408 217
rect 1442 183 1464 217
rect 1386 0 1464 183
rect 1494 217 1572 400
rect 1494 183 1516 217
rect 1550 183 1572 217
rect 1494 0 1572 183
rect 1602 217 1680 400
rect 1602 183 1624 217
rect 1658 183 1680 217
rect 1602 0 1680 183
rect 1710 217 1788 400
rect 1710 183 1732 217
rect 1766 183 1788 217
rect 1710 0 1788 183
rect 1818 217 1896 400
rect 1818 183 1840 217
rect 1874 183 1896 217
rect 1818 0 1896 183
rect 1926 217 2004 400
rect 1926 183 1948 217
rect 1982 183 2004 217
rect 1926 0 2004 183
rect 2034 217 2112 400
rect 2034 183 2056 217
rect 2090 183 2112 217
rect 2034 0 2112 183
rect 2142 217 2220 400
rect 2142 183 2164 217
rect 2198 183 2220 217
rect 2142 0 2220 183
rect 2250 217 2328 400
rect 2250 183 2272 217
rect 2306 183 2328 217
rect 2250 0 2328 183
rect 2358 217 2436 400
rect 2358 183 2380 217
rect 2414 183 2436 217
rect 2358 0 2436 183
rect 2466 217 2544 400
rect 2466 183 2488 217
rect 2522 183 2544 217
rect 2466 0 2544 183
rect 2574 217 2652 400
rect 2574 183 2596 217
rect 2630 183 2652 217
rect 2574 0 2652 183
rect 2682 217 2760 400
rect 2682 183 2704 217
rect 2738 183 2760 217
rect 2682 0 2760 183
rect 2790 217 2868 400
rect 2790 183 2812 217
rect 2846 183 2868 217
rect 2790 0 2868 183
rect 2898 217 2976 400
rect 2898 183 2920 217
rect 2954 183 2976 217
rect 2898 0 2976 183
rect 3006 217 3084 400
rect 3006 183 3028 217
rect 3062 183 3084 217
rect 3006 0 3084 183
rect 3114 217 3192 400
rect 3114 183 3136 217
rect 3170 183 3192 217
rect 3114 0 3192 183
rect 3222 217 3300 400
rect 3222 183 3244 217
rect 3278 183 3300 217
rect 3222 0 3300 183
rect 3330 217 3408 400
rect 3330 183 3352 217
rect 3386 183 3408 217
rect 3330 0 3408 183
rect 3438 217 3516 400
rect 3438 183 3460 217
rect 3494 183 3516 217
rect 3438 0 3516 183
rect 3546 217 3624 400
rect 3546 183 3568 217
rect 3602 183 3624 217
rect 3546 0 3624 183
rect 3654 217 3732 400
rect 3654 183 3676 217
rect 3710 183 3732 217
rect 3654 0 3732 183
rect 3762 217 3840 400
rect 3762 183 3784 217
rect 3818 183 3840 217
rect 3762 0 3840 183
rect 3870 217 3948 400
rect 3870 183 3892 217
rect 3926 183 3948 217
rect 3870 0 3948 183
rect 3978 217 4056 400
rect 3978 183 4000 217
rect 4034 183 4056 217
rect 3978 0 4056 183
rect 4086 217 4164 400
rect 4086 183 4108 217
rect 4142 183 4164 217
rect 4086 0 4164 183
rect 4194 217 4272 400
rect 4194 183 4216 217
rect 4250 183 4272 217
rect 4194 0 4272 183
rect 4302 217 4380 400
rect 4302 183 4324 217
rect 4358 183 4380 217
rect 4302 0 4380 183
rect 4410 217 4488 400
rect 4410 183 4432 217
rect 4466 183 4488 217
rect 4410 0 4488 183
rect 4518 217 4578 400
rect 4518 183 4536 217
rect 4570 183 4578 217
rect 4518 0 4578 183
<< pdiffc >>
rect 8 183 42 217
rect 112 183 146 217
rect 220 183 254 217
rect 328 183 362 217
rect 436 183 470 217
rect 544 183 578 217
rect 652 183 686 217
rect 760 183 794 217
rect 868 183 902 217
rect 976 183 1010 217
rect 1084 183 1118 217
rect 1192 183 1226 217
rect 1300 183 1334 217
rect 1408 183 1442 217
rect 1516 183 1550 217
rect 1624 183 1658 217
rect 1732 183 1766 217
rect 1840 183 1874 217
rect 1948 183 1982 217
rect 2056 183 2090 217
rect 2164 183 2198 217
rect 2272 183 2306 217
rect 2380 183 2414 217
rect 2488 183 2522 217
rect 2596 183 2630 217
rect 2704 183 2738 217
rect 2812 183 2846 217
rect 2920 183 2954 217
rect 3028 183 3062 217
rect 3136 183 3170 217
rect 3244 183 3278 217
rect 3352 183 3386 217
rect 3460 183 3494 217
rect 3568 183 3602 217
rect 3676 183 3710 217
rect 3784 183 3818 217
rect 3892 183 3926 217
rect 4000 183 4034 217
rect 4108 183 4142 217
rect 4216 183 4250 217
rect 4324 183 4358 217
rect 4432 183 4466 217
rect 4536 183 4570 217
<< poly >>
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 384 400 414 426
rect 492 400 522 426
rect 600 400 630 426
rect 708 400 738 426
rect 816 400 846 426
rect 924 400 954 426
rect 1032 400 1062 426
rect 1140 400 1170 426
rect 1248 400 1278 426
rect 1356 400 1386 426
rect 1464 400 1494 426
rect 1572 400 1602 426
rect 1680 400 1710 426
rect 1788 400 1818 426
rect 1896 400 1926 426
rect 2004 400 2034 426
rect 2112 400 2142 426
rect 2220 400 2250 426
rect 2328 400 2358 426
rect 2436 400 2466 426
rect 2544 400 2574 426
rect 2652 400 2682 426
rect 2760 400 2790 426
rect 2868 400 2898 426
rect 2976 400 3006 426
rect 3084 400 3114 426
rect 3192 400 3222 426
rect 3300 400 3330 426
rect 3408 400 3438 426
rect 3516 400 3546 426
rect 3624 400 3654 426
rect 3732 400 3762 426
rect 3840 400 3870 426
rect 3948 400 3978 426
rect 4056 400 4086 426
rect 4164 400 4194 426
rect 4272 400 4302 426
rect 4380 400 4410 426
rect 4488 400 4518 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 2328 -26 2358 0
rect 2436 -26 2466 0
rect 2544 -26 2574 0
rect 2652 -26 2682 0
rect 2760 -26 2790 0
rect 2868 -26 2898 0
rect 2976 -26 3006 0
rect 3084 -26 3114 0
rect 3192 -26 3222 0
rect 3300 -26 3330 0
rect 3408 -26 3438 0
rect 3516 -26 3546 0
rect 3624 -26 3654 0
rect 3732 -26 3762 0
rect 3840 -26 3870 0
rect 3948 -26 3978 0
rect 4056 -26 4086 0
rect 4164 -26 4194 0
rect 4272 -26 4302 0
rect 4380 -26 4410 0
rect 4488 -26 4518 0
rect 60 -56 4518 -26
<< locali >>
rect 8 217 42 233
rect 8 167 42 183
rect 112 217 146 233
rect 112 133 146 183
rect 220 217 254 233
rect 220 167 254 183
rect 328 217 362 233
rect 328 133 362 183
rect 436 217 470 233
rect 436 167 470 183
rect 544 217 578 233
rect 544 133 578 183
rect 652 217 686 233
rect 652 167 686 183
rect 760 217 794 233
rect 760 133 794 183
rect 868 217 902 233
rect 868 167 902 183
rect 976 217 1010 233
rect 976 133 1010 183
rect 1084 217 1118 233
rect 1084 167 1118 183
rect 1192 217 1226 233
rect 1192 133 1226 183
rect 1300 217 1334 233
rect 1300 167 1334 183
rect 1408 217 1442 233
rect 1408 133 1442 183
rect 1516 217 1550 233
rect 1516 167 1550 183
rect 1624 217 1658 233
rect 1624 133 1658 183
rect 1732 217 1766 233
rect 1732 167 1766 183
rect 1840 217 1874 233
rect 1840 133 1874 183
rect 1948 217 1982 233
rect 1948 167 1982 183
rect 2056 217 2090 233
rect 2056 133 2090 183
rect 2164 217 2198 233
rect 2164 167 2198 183
rect 2272 217 2306 233
rect 2272 133 2306 183
rect 2380 217 2414 233
rect 2380 167 2414 183
rect 2488 217 2522 233
rect 2488 133 2522 183
rect 2596 217 2630 233
rect 2596 167 2630 183
rect 2704 217 2738 233
rect 2704 133 2738 183
rect 2812 217 2846 233
rect 2812 167 2846 183
rect 2920 217 2954 233
rect 2920 133 2954 183
rect 3028 217 3062 233
rect 3028 167 3062 183
rect 3136 217 3170 233
rect 3136 133 3170 183
rect 3244 217 3278 233
rect 3244 167 3278 183
rect 3352 217 3386 233
rect 3352 133 3386 183
rect 3460 217 3494 233
rect 3460 167 3494 183
rect 3568 217 3602 233
rect 3568 133 3602 183
rect 3676 217 3710 233
rect 3676 167 3710 183
rect 3784 217 3818 233
rect 3784 133 3818 183
rect 3892 217 3926 233
rect 3892 167 3926 183
rect 4000 217 4034 233
rect 4000 133 4034 183
rect 4108 217 4142 233
rect 4108 167 4142 183
rect 4216 217 4250 233
rect 4216 133 4250 183
rect 4324 217 4358 233
rect 4324 167 4358 183
rect 4432 217 4466 233
rect 4432 133 4466 183
rect 4536 217 4570 233
rect 4536 167 4570 183
rect 112 99 4466 133
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_0
timestamp 1676037725
transform 1 0 4528 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_1
timestamp 1676037725
transform 1 0 4424 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_2
timestamp 1676037725
transform 1 0 4316 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_3
timestamp 1676037725
transform 1 0 4208 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_4
timestamp 1676037725
transform 1 0 4100 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_5
timestamp 1676037725
transform 1 0 3992 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_6
timestamp 1676037725
transform 1 0 3884 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_7
timestamp 1676037725
transform 1 0 3776 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_8
timestamp 1676037725
transform 1 0 3668 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_9
timestamp 1676037725
transform 1 0 3560 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_10
timestamp 1676037725
transform 1 0 3452 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_11
timestamp 1676037725
transform 1 0 3344 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_12
timestamp 1676037725
transform 1 0 3236 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_13
timestamp 1676037725
transform 1 0 3128 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_14
timestamp 1676037725
transform 1 0 3020 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_15
timestamp 1676037725
transform 1 0 2912 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_16
timestamp 1676037725
transform 1 0 2804 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_17
timestamp 1676037725
transform 1 0 2696 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_18
timestamp 1676037725
transform 1 0 2588 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_19
timestamp 1676037725
transform 1 0 2480 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_20
timestamp 1676037725
transform 1 0 2372 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_21
timestamp 1676037725
transform 1 0 2264 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_22
timestamp 1676037725
transform 1 0 2156 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_23
timestamp 1676037725
transform 1 0 2048 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_24
timestamp 1676037725
transform 1 0 1940 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_25
timestamp 1676037725
transform 1 0 1832 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_26
timestamp 1676037725
transform 1 0 1724 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_27
timestamp 1676037725
transform 1 0 1616 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_28
timestamp 1676037725
transform 1 0 1508 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_29
timestamp 1676037725
transform 1 0 1400 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_30
timestamp 1676037725
transform 1 0 1292 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_31
timestamp 1676037725
transform 1 0 1184 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_32
timestamp 1676037725
transform 1 0 1076 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_33
timestamp 1676037725
transform 1 0 968 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_34
timestamp 1676037725
transform 1 0 860 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_35
timestamp 1676037725
transform 1 0 752 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_36
timestamp 1676037725
transform 1 0 644 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_37
timestamp 1676037725
transform 1 0 536 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_38
timestamp 1676037725
transform 1 0 428 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_39
timestamp 1676037725
transform 1 0 320 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_40
timestamp 1676037725
transform 1 0 212 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_41
timestamp 1676037725
transform 1 0 104 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_42
timestamp 1676037725
transform 1 0 0 0 1 167
box 0 0 1 1
<< labels >>
rlabel locali s 1317 200 1317 200 4 S
rlabel locali s 237 200 237 200 4 S
rlabel locali s 3909 200 3909 200 4 S
rlabel locali s 3477 200 3477 200 4 S
rlabel locali s 4125 200 4125 200 4 S
rlabel locali s 1749 200 1749 200 4 S
rlabel locali s 4341 200 4341 200 4 S
rlabel locali s 4553 200 4553 200 4 S
rlabel locali s 2397 200 2397 200 4 S
rlabel locali s 453 200 453 200 4 S
rlabel locali s 2829 200 2829 200 4 S
rlabel locali s 885 200 885 200 4 S
rlabel locali s 1533 200 1533 200 4 S
rlabel locali s 3045 200 3045 200 4 S
rlabel locali s 2181 200 2181 200 4 S
rlabel locali s 1965 200 1965 200 4 S
rlabel locali s 2613 200 2613 200 4 S
rlabel locali s 1101 200 1101 200 4 S
rlabel locali s 669 200 669 200 4 S
rlabel locali s 25 200 25 200 4 S
rlabel locali s 3693 200 3693 200 4 S
rlabel locali s 3261 200 3261 200 4 S
rlabel locali s 2289 116 2289 116 4 D
rlabel poly s 2289 -41 2289 -41 4 G
<< properties >>
string FIXED_BBOX -54 -56 4632 116
string GDS_END 149956
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 139826
<< end >>
