magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 365 157 551 203
rect 1 21 551 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 267 47 297 131
rect 345 47 375 131
rect 443 47 473 177
<< scpmoshvt >>
rect 79 413 109 497
rect 177 413 207 497
rect 265 413 295 497
rect 443 297 473 497
<< ndiff >>
rect 391 131 443 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 106 161 131
rect 109 72 119 106
rect 153 72 161 106
rect 109 47 161 72
rect 215 106 267 131
rect 215 72 223 106
rect 257 72 267 106
rect 215 47 267 72
rect 297 47 345 131
rect 375 111 443 131
rect 375 77 399 111
rect 433 77 443 111
rect 375 47 443 77
rect 473 127 525 177
rect 473 93 483 127
rect 517 93 525 127
rect 473 47 525 93
<< pdiff >>
rect 27 462 79 497
rect 27 428 35 462
rect 69 428 79 462
rect 27 413 79 428
rect 109 471 177 497
rect 109 437 119 471
rect 153 437 177 471
rect 109 413 177 437
rect 207 462 265 497
rect 207 428 219 462
rect 253 428 265 462
rect 207 413 265 428
rect 295 483 443 497
rect 295 449 315 483
rect 349 449 383 483
rect 417 449 443 483
rect 295 413 443 449
rect 393 297 443 413
rect 473 457 525 497
rect 473 423 483 457
rect 517 423 525 457
rect 473 384 525 423
rect 473 350 483 384
rect 517 350 525 384
rect 473 297 525 350
<< ndiffc >>
rect 35 72 69 106
rect 119 72 153 106
rect 223 72 257 106
rect 399 77 433 111
rect 483 93 517 127
<< pdiffc >>
rect 35 428 69 462
rect 119 437 153 471
rect 219 428 253 462
rect 315 449 349 483
rect 383 449 417 483
rect 483 423 517 457
rect 483 350 517 384
<< poly >>
rect 79 497 109 523
rect 177 497 207 523
rect 265 497 295 523
rect 443 497 473 523
rect 79 265 109 413
rect 39 249 109 265
rect 39 215 55 249
rect 89 215 109 249
rect 39 199 109 215
rect 79 131 109 199
rect 177 227 207 413
rect 265 379 295 413
rect 265 363 363 379
rect 265 329 312 363
rect 346 329 363 363
rect 265 305 363 329
rect 289 282 363 305
rect 289 233 375 282
rect 443 265 473 297
rect 177 211 246 227
rect 177 177 196 211
rect 230 191 246 211
rect 230 177 297 191
rect 177 161 297 177
rect 267 131 297 161
rect 345 131 375 233
rect 417 249 473 265
rect 417 215 427 249
rect 461 215 473 249
rect 417 197 473 215
rect 443 177 473 197
rect 79 21 109 47
rect 267 21 297 47
rect 345 21 375 47
rect 443 21 473 47
<< polycont >>
rect 55 215 89 249
rect 312 329 346 363
rect 196 177 230 211
rect 427 215 461 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 35 462 69 489
rect 103 471 169 527
rect 103 437 119 471
rect 153 437 169 471
rect 204 462 261 484
rect 35 403 69 428
rect 204 428 219 462
rect 253 428 261 462
rect 297 483 434 527
rect 297 449 315 483
rect 349 449 383 483
rect 417 449 434 483
rect 297 433 434 449
rect 470 457 531 473
rect 35 357 170 403
rect 29 249 89 323
rect 29 215 55 249
rect 29 153 89 215
rect 123 227 170 357
rect 204 295 261 428
rect 470 423 483 457
rect 517 423 531 457
rect 296 363 435 391
rect 296 329 312 363
rect 346 329 435 363
rect 470 384 531 423
rect 470 350 483 384
rect 517 350 531 384
rect 470 316 531 350
rect 204 265 376 295
rect 204 261 461 265
rect 264 249 461 261
rect 123 211 230 227
rect 123 177 196 211
rect 123 161 230 177
rect 264 215 427 249
rect 264 189 461 215
rect 123 131 167 161
rect 18 106 85 118
rect 18 72 35 106
rect 69 72 85 106
rect 18 17 85 72
rect 119 106 167 131
rect 264 122 298 189
rect 496 155 531 316
rect 153 72 167 106
rect 119 56 167 72
rect 223 106 298 122
rect 483 127 531 155
rect 257 83 298 106
rect 370 111 449 116
rect 223 54 257 72
rect 370 77 399 111
rect 433 77 449 111
rect 370 17 449 77
rect 517 93 531 127
rect 483 51 531 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 489 357 523 391 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 305 357 339 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 489 85 523 119 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 397 357 431 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 489 425 523 459 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and2b_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 3852686
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3847210
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 13.800 13.600 
<< end >>
