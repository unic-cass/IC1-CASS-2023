magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 98 157 459 203
rect 1 21 459 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 256 47 286 177
rect 351 47 381 177
<< scpmoshvt >>
rect 79 369 109 497
rect 174 297 204 497
rect 351 297 381 497
<< ndiff >>
rect 124 131 256 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 256 131
rect 109 55 131 89
rect 165 55 199 89
rect 233 55 256 89
rect 109 47 256 55
rect 286 47 351 177
rect 381 103 433 177
rect 381 69 391 103
rect 425 69 433 103
rect 381 47 433 69
<< pdiff >>
rect 27 450 79 497
rect 27 416 35 450
rect 69 416 79 450
rect 27 369 79 416
rect 109 489 174 497
rect 109 455 124 489
rect 158 455 174 489
rect 109 369 174 455
rect 124 297 174 369
rect 204 297 351 497
rect 381 477 433 497
rect 381 443 391 477
rect 425 443 433 477
rect 381 409 433 443
rect 381 375 391 409
rect 425 375 433 409
rect 381 297 433 375
<< ndiffc >>
rect 35 72 69 106
rect 131 55 165 89
rect 199 55 233 89
rect 391 69 425 103
<< pdiffc >>
rect 35 416 69 450
rect 124 455 158 489
rect 391 443 425 477
rect 391 375 425 409
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 351 497 381 523
rect 79 282 109 369
rect 174 282 204 297
rect 79 265 204 282
rect 351 265 381 297
rect 54 252 204 265
rect 54 249 109 252
rect 54 215 64 249
rect 98 215 109 249
rect 54 199 109 215
rect 246 249 309 265
rect 246 215 256 249
rect 290 215 309 249
rect 246 199 309 215
rect 351 249 438 265
rect 351 215 394 249
rect 428 215 438 249
rect 351 199 438 215
rect 79 131 109 199
rect 256 177 286 199
rect 351 177 381 199
rect 79 21 109 47
rect 256 21 286 47
rect 351 21 381 47
<< polycont >>
rect 64 215 98 249
rect 256 215 290 249
rect 394 215 428 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 450 74 493
rect 17 416 35 450
rect 69 416 74 450
rect 108 489 174 527
rect 108 455 124 489
rect 158 455 174 489
rect 108 447 174 455
rect 208 477 443 493
rect 17 413 74 416
rect 208 443 391 477
rect 425 443 443 477
rect 17 379 174 413
rect 17 249 102 345
rect 17 215 64 249
rect 98 215 102 249
rect 17 191 102 215
rect 137 323 174 379
rect 208 409 443 443
rect 208 375 391 409
rect 425 375 443 409
rect 208 357 443 375
rect 137 249 290 323
rect 137 215 256 249
rect 137 157 290 215
rect 17 123 290 157
rect 17 106 74 123
rect 17 72 35 106
rect 69 72 74 106
rect 324 119 360 357
rect 394 249 443 323
rect 428 215 443 249
rect 394 153 443 215
rect 324 103 443 119
rect 17 51 74 72
rect 108 55 131 89
rect 165 55 199 89
rect 233 55 288 89
rect 108 17 288 55
rect 324 69 391 103
rect 425 69 443 103
rect 324 51 443 69
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 212 357 246 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 212 425 246 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 304 357 338 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 304 425 338 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 396 425 430 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 396 357 430 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 396 85 430 119 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 396 153 430 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 396 221 430 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 396 289 430 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 einvn_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 2965730
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2960664
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
