magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -66 377 1986 897
<< pwell >>
rect 1650 217 1916 283
rect 6 43 1916 217
rect -26 -43 1946 43
<< locali >>
rect 114 386 180 520
rect 121 235 359 280
rect 1747 435 1895 751
rect 1503 356 1569 371
rect 1503 162 1624 356
rect 1828 99 1895 435
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 114 735 304 741
rect 28 350 78 722
rect 114 701 120 735
rect 154 701 192 735
rect 226 701 264 735
rect 298 701 304 735
rect 560 735 750 741
rect 114 556 304 701
rect 340 439 406 722
rect 560 701 566 735
rect 600 701 638 735
rect 672 701 710 735
rect 744 701 750 735
rect 458 509 524 649
rect 560 545 750 701
rect 1141 735 1331 741
rect 1141 701 1147 735
rect 1181 701 1219 735
rect 1253 701 1291 735
rect 1325 701 1331 735
rect 912 579 978 649
rect 912 545 1105 579
rect 458 475 957 509
rect 923 459 957 475
rect 340 405 887 439
rect 325 350 731 369
rect 28 335 731 350
rect 28 316 359 335
rect 767 321 887 405
rect 923 393 1035 459
rect 28 99 78 316
rect 767 299 801 321
rect 395 265 801 299
rect 923 279 957 393
rect 395 199 429 265
rect 837 245 957 279
rect 1071 269 1105 545
rect 1141 451 1331 701
rect 1514 735 1704 751
rect 1514 701 1520 735
rect 1554 701 1592 735
rect 1626 701 1664 735
rect 1698 701 1704 735
rect 1392 441 1478 601
rect 1514 477 1704 701
rect 1392 415 1694 441
rect 1162 407 1694 415
rect 1162 381 1426 407
rect 1162 305 1228 381
rect 1290 269 1356 345
rect 837 229 899 245
rect 114 113 304 199
rect 114 79 120 113
rect 154 79 192 113
rect 226 79 264 113
rect 298 79 304 113
rect 340 99 429 199
rect 474 195 899 229
rect 993 235 1356 269
rect 993 199 1027 235
rect 1392 199 1426 381
rect 1660 399 1694 407
rect 474 99 524 195
rect 560 113 750 159
rect 114 73 304 79
rect 560 79 566 113
rect 600 79 638 113
rect 672 79 710 113
rect 744 79 750 113
rect 935 99 1027 199
rect 1109 113 1299 199
rect 560 73 750 79
rect 1109 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1259 113
rect 1293 79 1299 113
rect 1351 99 1426 199
rect 1660 333 1726 399
rect 1660 113 1778 265
rect 1109 73 1299 79
rect 1660 79 1666 113
rect 1700 79 1738 113
rect 1772 79 1778 113
rect 1660 73 1778 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 120 701 154 735
rect 192 701 226 735
rect 264 701 298 735
rect 566 701 600 735
rect 638 701 672 735
rect 710 701 744 735
rect 1147 701 1181 735
rect 1219 701 1253 735
rect 1291 701 1325 735
rect 1520 701 1554 735
rect 1592 701 1626 735
rect 1664 701 1698 735
rect 120 79 154 113
rect 192 79 226 113
rect 264 79 298 113
rect 566 79 600 113
rect 638 79 672 113
rect 710 79 744 113
rect 1115 79 1149 113
rect 1187 79 1221 113
rect 1259 79 1293 113
rect 1666 79 1700 113
rect 1738 79 1772 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 831 1920 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 0 791 1920 797
rect 0 735 1920 763
rect 0 701 120 735
rect 154 701 192 735
rect 226 701 264 735
rect 298 701 566 735
rect 600 701 638 735
rect 672 701 710 735
rect 744 701 1147 735
rect 1181 701 1219 735
rect 1253 701 1291 735
rect 1325 701 1520 735
rect 1554 701 1592 735
rect 1626 701 1664 735
rect 1698 701 1920 735
rect 0 689 1920 701
rect 0 113 1920 125
rect 0 79 120 113
rect 154 79 192 113
rect 226 79 264 113
rect 298 79 566 113
rect 600 79 638 113
rect 672 79 710 113
rect 744 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1259 113
rect 1293 79 1666 113
rect 1700 79 1738 113
rect 1772 79 1920 113
rect 0 51 1920 79
rect 0 17 1920 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -23 1920 -17
<< labels >>
rlabel locali s 114 386 180 520 6 D
port 1 nsew signal input
rlabel locali s 121 235 359 280 6 GATE
port 2 nsew clock input
rlabel locali s 1503 162 1624 356 6 RESET_B
port 3 nsew signal input
rlabel locali s 1503 356 1569 371 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 51 1920 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 1920 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 1946 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 6 43 1916 217 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1650 217 1916 283 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 1920 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 1986 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 1920 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 1828 99 1895 435 6 Q
port 8 nsew signal output
rlabel locali s 1747 435 1895 751 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1920 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1203658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1183922
<< end >>
